module intadder_35_freq500_uid41
  (input  clk,
   input  [34:0] x,
   input  [34:0] y,
   input  cin,
   output [34:0] r);
  wire [34:0] rtmp;
  wire cin_d1;
  wire [34:0] n4763;
  wire [34:0] n4764;
  wire [34:0] n4765;
  reg n4766;
  assign r = rtmp; //(module output)
  /* fplog32.vhdl:1947:8  */
  assign rtmp = n4765; // (signal)
  /* fplog32.vhdl:1949:8  */
  assign cin_d1 = n4766; // (signal)
  /* fplog32.vhdl:1958:14  */
  assign n4763 = x + y;
  /* fplog32.vhdl:1958:18  */
  assign n4764 = {34'b0, cin_d1};  //  uext
  /* fplog32.vhdl:1958:18  */
  assign n4765 = n4763 + n4764;
  /* fplog32.vhdl:1954:10  */
  always @(posedge clk)
    n4766 <= cin;
endmodule

module fixrealkcm_freq500_uid31_t1_freq500_uid37
  (input  [2:0] x,
   output [29:0] y);
  wire [29:0] y0;
  wire [29:0] y1;
  wire n4732;
  wire n4735;
  wire n4738;
  wire n4741;
  wire n4744;
  wire n4747;
  wire n4750;
  wire n4753;
  wire [7:0] n4755;
  reg [29:0] n4756;
  assign y = y1; //(module output)
  /* fplog32.vhdl:822:8  */
  assign y0 = n4756; // (signal)
  /* fplog32.vhdl:824:8  */
  assign y1 = y0; // (signal)
  /* fplog32.vhdl:828:40  */
  assign n4732 = x == 3'b000;
  /* fplog32.vhdl:829:40  */
  assign n4735 = x == 3'b001;
  /* fplog32.vhdl:830:40  */
  assign n4738 = x == 3'b010;
  /* fplog32.vhdl:831:40  */
  assign n4741 = x == 3'b011;
  /* fplog32.vhdl:832:40  */
  assign n4744 = x == 3'b100;
  /* fplog32.vhdl:833:40  */
  assign n4747 = x == 3'b101;
  /* fplog32.vhdl:834:40  */
  assign n4750 = x == 3'b110;
  /* fplog32.vhdl:835:40  */
  assign n4753 = x == 3'b111;
  assign n4755 = {n4753, n4750, n4747, n4744, n4741, n4738, n4735, n4732};
  /* fplog32.vhdl:827:4  */
  always @*
    case (n4755)
      8'b10000000: n4756 = 30'b100110110100001111010100111110;
      8'b01000000: n4756 = 30'b100001010001010110010001111110;
      8'b00100000: n4756 = 30'b011011101110011101001110111111;
      8'b00010000: n4756 = 30'b010110001011100100001011111111;
      8'b00001000: n4756 = 30'b010000101000101011001000111111;
      8'b00000100: n4756 = 30'b001011000101110010000101111111;
      8'b00000010: n4756 = 30'b000101100010111001000011000000;
      8'b00000001: n4756 = 30'b000000000000000000000000000000;
      default: n4756 = 30'bX;
    endcase
endmodule

module fixrealkcm_freq500_uid31_t0_freq500_uid34
  (input  [4:0] x,
   output [34:0] y);
  wire [34:0] y0;
  wire [34:0] y1;
  wire n4632;
  wire n4635;
  wire n4638;
  wire n4641;
  wire n4644;
  wire n4647;
  wire n4650;
  wire n4653;
  wire n4656;
  wire n4659;
  wire n4662;
  wire n4665;
  wire n4668;
  wire n4671;
  wire n4674;
  wire n4677;
  wire n4680;
  wire n4683;
  wire n4686;
  wire n4689;
  wire n4692;
  wire n4695;
  wire n4698;
  wire n4701;
  wire n4704;
  wire n4707;
  wire n4710;
  wire n4713;
  wire n4716;
  wire n4719;
  wire n4722;
  wire n4725;
  wire [31:0] n4727;
  reg [34:0] n4728;
  assign y = y1; //(module output)
  /* fplog32.vhdl:750:8  */
  assign y0 = n4728; // (signal)
  /* fplog32.vhdl:752:8  */
  assign y1 = y0; // (signal)
  /* fplog32.vhdl:756:45  */
  assign n4632 = x == 5'b00000;
  /* fplog32.vhdl:757:45  */
  assign n4635 = x == 5'b00001;
  /* fplog32.vhdl:758:45  */
  assign n4638 = x == 5'b00010;
  /* fplog32.vhdl:759:45  */
  assign n4641 = x == 5'b00011;
  /* fplog32.vhdl:760:45  */
  assign n4644 = x == 5'b00100;
  /* fplog32.vhdl:761:45  */
  assign n4647 = x == 5'b00101;
  /* fplog32.vhdl:762:45  */
  assign n4650 = x == 5'b00110;
  /* fplog32.vhdl:763:45  */
  assign n4653 = x == 5'b00111;
  /* fplog32.vhdl:764:45  */
  assign n4656 = x == 5'b01000;
  /* fplog32.vhdl:765:45  */
  assign n4659 = x == 5'b01001;
  /* fplog32.vhdl:766:45  */
  assign n4662 = x == 5'b01010;
  /* fplog32.vhdl:767:45  */
  assign n4665 = x == 5'b01011;
  /* fplog32.vhdl:768:45  */
  assign n4668 = x == 5'b01100;
  /* fplog32.vhdl:769:45  */
  assign n4671 = x == 5'b01101;
  /* fplog32.vhdl:770:45  */
  assign n4674 = x == 5'b01110;
  /* fplog32.vhdl:771:45  */
  assign n4677 = x == 5'b01111;
  /* fplog32.vhdl:772:45  */
  assign n4680 = x == 5'b10000;
  /* fplog32.vhdl:773:45  */
  assign n4683 = x == 5'b10001;
  /* fplog32.vhdl:774:45  */
  assign n4686 = x == 5'b10010;
  /* fplog32.vhdl:775:45  */
  assign n4689 = x == 5'b10011;
  /* fplog32.vhdl:776:45  */
  assign n4692 = x == 5'b10100;
  /* fplog32.vhdl:777:45  */
  assign n4695 = x == 5'b10101;
  /* fplog32.vhdl:778:45  */
  assign n4698 = x == 5'b10110;
  /* fplog32.vhdl:779:45  */
  assign n4701 = x == 5'b10111;
  /* fplog32.vhdl:780:45  */
  assign n4704 = x == 5'b11000;
  /* fplog32.vhdl:781:45  */
  assign n4707 = x == 5'b11001;
  /* fplog32.vhdl:782:45  */
  assign n4710 = x == 5'b11010;
  /* fplog32.vhdl:783:45  */
  assign n4713 = x == 5'b11011;
  /* fplog32.vhdl:784:45  */
  assign n4716 = x == 5'b11100;
  /* fplog32.vhdl:785:45  */
  assign n4719 = x == 5'b11101;
  /* fplog32.vhdl:786:45  */
  assign n4722 = x == 5'b11110;
  /* fplog32.vhdl:787:45  */
  assign n4725 = x == 5'b11111;
  assign n4727 = {n4725, n4722, n4719, n4716, n4713, n4710, n4707, n4704, n4701, n4698, n4695, n4692, n4689, n4686, n4683, n4680, n4677, n4674, n4671, n4668, n4665, n4662, n4659, n4656, n4653, n4650, n4647, n4644, n4641, n4638, n4635, n4632};
  /* fplog32.vhdl:755:4  */
  always @*
    case (n4727)
      32'b10000000000000000000000000000000: n4728 = 35'b10101011111001101000011100111000001;
      32'b01000000000000000000000000000000: n4728 = 35'b10100110010110101111011001111000011;
      32'b00100000000000000000000000000000: n4728 = 35'b10100000110011110110010110111000101;
      32'b00010000000000000000000000000000: n4728 = 35'b10011011010000111101010011111000111;
      32'b00001000000000000000000000000000: n4728 = 35'b10010101101110000100010000111001001;
      32'b00000100000000000000000000000000: n4728 = 35'b10010000001011001011001101111001011;
      32'b00000010000000000000000000000000: n4728 = 35'b10001010101000010010001010111001101;
      32'b00000001000000000000000000000000: n4728 = 35'b10000101000101011001000111111001111;
      32'b00000000100000000000000000000000: n4728 = 35'b01111111100010100000000100111010001;
      32'b00000000010000000000000000000000: n4728 = 35'b01111001111111100111000001111010011;
      32'b00000000001000000000000000000000: n4728 = 35'b01110100011100101101111110111010101;
      32'b00000000000100000000000000000000: n4728 = 35'b01101110111001110100111011111010111;
      32'b00000000000010000000000000000000: n4728 = 35'b01101001010110111011111000111011001;
      32'b00000000000001000000000000000000: n4728 = 35'b01100011110100000010110101111011011;
      32'b00000000000000100000000000000000: n4728 = 35'b01011110010001001001110010111011101;
      32'b00000000000000010000000000000000: n4728 = 35'b01011000101110010000101111111011111;
      32'b00000000000000001000000000000000: n4728 = 35'b01010011001011010111101100111100001;
      32'b00000000000000000100000000000000: n4728 = 35'b01001101101000011110101001111100011;
      32'b00000000000000000010000000000000: n4728 = 35'b01001000000101100101100110111100101;
      32'b00000000000000000001000000000000: n4728 = 35'b01000010100010101100100011111100111;
      32'b00000000000000000000100000000000: n4728 = 35'b00111100111111110011100000111101010;
      32'b00000000000000000000010000000000: n4728 = 35'b00110111011100111010011101111101100;
      32'b00000000000000000000001000000000: n4728 = 35'b00110001111010000001011010111101110;
      32'b00000000000000000000000100000000: n4728 = 35'b00101100010111001000010111111110000;
      32'b00000000000000000000000010000000: n4728 = 35'b00100110110100001111010100111110010;
      32'b00000000000000000000000001000000: n4728 = 35'b00100001010001010110010001111110100;
      32'b00000000000000000000000000100000: n4728 = 35'b00011011101110011101001110111110110;
      32'b00000000000000000000000000010000: n4728 = 35'b00010110001011100100001011111111000;
      32'b00000000000000000000000000001000: n4728 = 35'b00010000101000101011001000111111010;
      32'b00000000000000000000000000000100: n4728 = 35'b00001011000101110010000101111111100;
      32'b00000000000000000000000000000010: n4728 = 35'b00000101100010111001000010111111110;
      32'b00000000000000000000000000000001: n4728 = 35'b00000000000000000000000000000000000;
      default: n4728 = 35'bX;
    endcase
endmodule

module intadder_31_freq500_uid52
  (input  clk,
   input  [30:0] x,
   input  [30:0] y,
   input  cin,
   output [30:0] r);
  wire cin_1;
  wire cin_1_d1;
  wire cin_1_d2;
  wire cin_1_d3;
  wire cin_1_d4;
  wire cin_1_d5;
  wire cin_1_d6;
  wire cin_1_d7;
  wire cin_1_d8;
  wire cin_1_d9;
  wire cin_1_d10;
  wire cin_1_d11;
  wire cin_1_d12;
  wire [31:0] x_1;
  wire [31:0] x_1_d1;
  wire [31:0] y_1;
  wire [31:0] y_1_d1;
  wire [31:0] s_1;
  wire [30:0] r_1;
  wire [31:0] n4608;
  wire [31:0] n4610;
  wire [31:0] n4611;
  wire [31:0] n4612;
  wire [31:0] n4613;
  wire [30:0] n4614;
  reg n4615;
  reg n4616;
  reg n4617;
  reg n4618;
  reg n4619;
  reg n4620;
  reg n4621;
  reg n4622;
  reg n4623;
  reg n4624;
  reg n4625;
  reg n4626;
  reg [31:0] n4627;
  reg [31:0] n4628;
  assign r = r_1; //(module output)
  /* fplog32.vhdl:2604:15  */
  assign cin_1_d1 = n4615; // (signal)
  /* fplog32.vhdl:2604:25  */
  assign cin_1_d2 = n4616; // (signal)
  /* fplog32.vhdl:2604:35  */
  assign cin_1_d3 = n4617; // (signal)
  /* fplog32.vhdl:2604:45  */
  assign cin_1_d4 = n4618; // (signal)
  /* fplog32.vhdl:2604:55  */
  assign cin_1_d5 = n4619; // (signal)
  /* fplog32.vhdl:2604:65  */
  assign cin_1_d6 = n4620; // (signal)
  /* fplog32.vhdl:2604:75  */
  assign cin_1_d7 = n4621; // (signal)
  /* fplog32.vhdl:2604:85  */
  assign cin_1_d8 = n4622; // (signal)
  /* fplog32.vhdl:2604:95  */
  assign cin_1_d9 = n4623; // (signal)
  /* fplog32.vhdl:2604:105  */
  assign cin_1_d10 = n4624; // (signal)
  /* fplog32.vhdl:2604:116  */
  assign cin_1_d11 = n4625; // (signal)
  /* fplog32.vhdl:2604:127  */
  assign cin_1_d12 = n4626; // (signal)
  /* fplog32.vhdl:2606:8  */
  assign x_1 = n4608; // (signal)
  /* fplog32.vhdl:2606:13  */
  assign x_1_d1 = n4627; // (signal)
  /* fplog32.vhdl:2608:8  */
  assign y_1 = n4610; // (signal)
  /* fplog32.vhdl:2608:13  */
  assign y_1_d1 = n4628; // (signal)
  /* fplog32.vhdl:2610:8  */
  assign s_1 = n4613; // (signal)
  /* fplog32.vhdl:2612:8  */
  assign r_1 = n4614; // (signal)
  /* fplog32.vhdl:2635:15  */
  assign n4608 = {1'b0, x};
  /* fplog32.vhdl:2636:15  */
  assign n4610 = {1'b0, y};
  /* fplog32.vhdl:2637:18  */
  assign n4611 = x_1_d1 + y_1_d1;
  /* fplog32.vhdl:2637:27  */
  assign n4612 = {31'b0, cin_1_d12};  //  uext
  /* fplog32.vhdl:2637:27  */
  assign n4613 = n4611 + n4612;
  /* fplog32.vhdl:2638:14  */
  assign n4614 = s_1[30:0]; // extract
  /* fplog32.vhdl:2617:10  */
  always @(posedge clk)
    n4615 <= cin_1;
  /* fplog32.vhdl:2617:10  */
  always @(posedge clk)
    n4616 <= cin_1_d1;
  /* fplog32.vhdl:2617:10  */
  always @(posedge clk)
    n4617 <= cin_1_d2;
  /* fplog32.vhdl:2617:10  */
  always @(posedge clk)
    n4618 <= cin_1_d3;
  /* fplog32.vhdl:2617:10  */
  always @(posedge clk)
    n4619 <= cin_1_d4;
  /* fplog32.vhdl:2617:10  */
  always @(posedge clk)
    n4620 <= cin_1_d5;
  /* fplog32.vhdl:2617:10  */
  always @(posedge clk)
    n4621 <= cin_1_d6;
  /* fplog32.vhdl:2617:10  */
  always @(posedge clk)
    n4622 <= cin_1_d7;
  /* fplog32.vhdl:2617:10  */
  always @(posedge clk)
    n4623 <= cin_1_d8;
  /* fplog32.vhdl:2617:10  */
  always @(posedge clk)
    n4624 <= cin_1_d9;
  /* fplog32.vhdl:2617:10  */
  always @(posedge clk)
    n4625 <= cin_1_d10;
  /* fplog32.vhdl:2617:10  */
  always @(posedge clk)
    n4626 <= cin_1_d11;
  /* fplog32.vhdl:2617:10  */
  always @(posedge clk)
    n4627 <= x_1;
  /* fplog32.vhdl:2617:10  */
  always @(posedge clk)
    n4628 <= y_1;
endmodule

module intadder_29_freq500_uid49
  (input  clk,
   input  [28:0] x,
   input  [28:0] y,
   input  cin,
   output [28:0] r);
  wire [28:0] rtmp;
  wire [28:0] x_d1;
  wire [28:0] x_d2;
  wire cin_d1;
  wire cin_d2;
  wire cin_d3;
  wire cin_d4;
  wire cin_d5;
  wire cin_d6;
  wire [28:0] n4577;
  wire [28:0] n4578;
  wire [28:0] n4579;
  reg [28:0] n4580;
  reg [28:0] n4581;
  reg n4582;
  reg n4583;
  reg n4584;
  reg n4585;
  reg n4586;
  reg n4587;
  assign r = rtmp; //(module output)
  /* fplog32.vhdl:2548:8  */
  assign rtmp = n4579; // (signal)
  /* fplog32.vhdl:2550:8  */
  assign x_d1 = n4580; // (signal)
  /* fplog32.vhdl:2550:14  */
  assign x_d2 = n4581; // (signal)
  /* fplog32.vhdl:2552:8  */
  assign cin_d1 = n4582; // (signal)
  /* fplog32.vhdl:2552:16  */
  assign cin_d2 = n4583; // (signal)
  /* fplog32.vhdl:2552:24  */
  assign cin_d3 = n4584; // (signal)
  /* fplog32.vhdl:2552:32  */
  assign cin_d4 = n4585; // (signal)
  /* fplog32.vhdl:2552:40  */
  assign cin_d5 = n4586; // (signal)
  /* fplog32.vhdl:2552:48  */
  assign cin_d6 = n4587; // (signal)
  /* fplog32.vhdl:2568:17  */
  assign n4577 = x_d2 + y;
  /* fplog32.vhdl:2568:21  */
  assign n4578 = {28'b0, cin_d6};  //  uext
  /* fplog32.vhdl:2568:21  */
  assign n4579 = n4577 + n4578;
  /* fplog32.vhdl:2557:10  */
  always @(posedge clk)
    n4580 <= x;
  /* fplog32.vhdl:2557:10  */
  always @(posedge clk)
    n4581 <= x_d1;
  /* fplog32.vhdl:2557:10  */
  always @(posedge clk)
    n4582 <= cin;
  /* fplog32.vhdl:2557:10  */
  always @(posedge clk)
    n4583 <= cin_d1;
  /* fplog32.vhdl:2557:10  */
  always @(posedge clk)
    n4584 <= cin_d2;
  /* fplog32.vhdl:2557:10  */
  always @(posedge clk)
    n4585 <= cin_d3;
  /* fplog32.vhdl:2557:10  */
  always @(posedge clk)
    n4586 <= cin_d4;
  /* fplog32.vhdl:2557:10  */
  always @(posedge clk)
    n4587 <= cin_d5;
endmodule

module rightshifter16_by_max_15_freq500_uid47
  (input  clk,
   input  [15:0] x,
   input  [3:0] s,
   output [30:0] r);
  wire [3:0] ps;
  wire [3:0] ps_d1;
  wire [3:0] ps_d2;
  wire [3:0] ps_d3;
  wire [15:0] level0;
  wire [16:0] level1;
  wire [18:0] level2;
  wire [22:0] level3;
  wire [22:0] level3_d1;
  wire [30:0] level4;
  wire [16:0] n4537;
  wire n4538;
  wire [16:0] n4539;
  wire [16:0] n4541;
  wire [18:0] n4543;
  wire n4544;
  wire [18:0] n4545;
  wire [18:0] n4547;
  wire [22:0] n4549;
  wire n4550;
  wire [22:0] n4551;
  wire [22:0] n4553;
  wire [30:0] n4555;
  wire n4556;
  wire [30:0] n4557;
  wire [30:0] n4559;
  reg [3:0] n4560;
  reg [3:0] n4561;
  reg [3:0] n4562;
  reg [22:0] n4563;
  assign r = level4; //(module output)
  /* fplog32.vhdl:2485:12  */
  assign ps_d1 = n4560; // (signal)
  /* fplog32.vhdl:2485:19  */
  assign ps_d2 = n4561; // (signal)
  /* fplog32.vhdl:2485:26  */
  assign ps_d3 = n4562; // (signal)
  /* fplog32.vhdl:2489:8  */
  assign level1 = n4539; // (signal)
  /* fplog32.vhdl:2491:8  */
  assign level2 = n4545; // (signal)
  /* fplog32.vhdl:2493:8  */
  assign level3 = n4551; // (signal)
  /* fplog32.vhdl:2493:16  */
  assign level3_d1 = n4563; // (signal)
  /* fplog32.vhdl:2495:8  */
  assign level4 = n4557; // (signal)
  /* fplog32.vhdl:2509:35  */
  assign n4537 = {1'b0, level0};
  /* fplog32.vhdl:2509:54  */
  assign n4538 = ps_d2[0]; // extract
  /* fplog32.vhdl:2509:44  */
  assign n4539 = n4538 ? n4537 : n4541;
  /* fplog32.vhdl:2509:79  */
  assign n4541 = {level0, 1'b0};
  /* fplog32.vhdl:2510:35  */
  assign n4543 = {2'b00, level1};
  /* fplog32.vhdl:2510:54  */
  assign n4544 = ps_d2[1]; // extract
  /* fplog32.vhdl:2510:44  */
  assign n4545 = n4544 ? n4543 : n4547;
  /* fplog32.vhdl:2510:79  */
  assign n4547 = {level1, 2'b00};
  /* fplog32.vhdl:2511:35  */
  assign n4549 = {4'b0000, level2};
  /* fplog32.vhdl:2511:54  */
  assign n4550 = ps_d2[2]; // extract
  /* fplog32.vhdl:2511:44  */
  assign n4551 = n4550 ? n4549 : n4553;
  /* fplog32.vhdl:2511:79  */
  assign n4553 = {level2, 4'b0000};
  /* fplog32.vhdl:2512:35  */
  assign n4555 = {8'b00000000, level3_d1};
  /* fplog32.vhdl:2512:57  */
  assign n4556 = ps_d3[3]; // extract
  /* fplog32.vhdl:2512:47  */
  assign n4557 = n4556 ? n4555 : n4559;
  /* fplog32.vhdl:2512:85  */
  assign n4559 = {level3_d1, 8'b00000000};
  /* fplog32.vhdl:2500:10  */
  always @(posedge clk)
    n4560 <= ps;
  /* fplog32.vhdl:2500:10  */
  always @(posedge clk)
    n4561 <= ps_d1;
  /* fplog32.vhdl:2500:10  */
  always @(posedge clk)
    n4562 <= ps_d2;
  /* fplog32.vhdl:2500:10  */
  always @(posedge clk)
    n4563 <= level3;
endmodule

module normalizer_z_48_40_19_freq500_uid45
  (input  clk,
   input  [47:0] x,
   output [4:0] count,
   output [39:0] r);
  wire [47:0] level5;
  wire [47:0] level5_d1;
  wire count4;
  wire count4_d1;
  wire count4_d2;
  wire [47:0] level4;
  wire [47:0] level4_d1;
  wire count3;
  wire count3_d1;
  wire count3_d2;
  wire [46:0] level3;
  wire count2;
  wire count2_d1;
  wire [42:0] level2;
  wire [42:0] level2_d1;
  wire count1;
  wire count1_d1;
  wire [40:0] level1;
  wire count0;
  wire [39:0] level0;
  wire [4:0] scount;
  wire [15:0] n4462;
  wire n4464;
  wire n4465;
  wire n4467;
  wire [47:0] n4468;
  wire [31:0] n4469;
  wire [47:0] n4471;
  wire [7:0] n4473;
  wire n4475;
  wire n4476;
  wire [46:0] n4478;
  wire n4479;
  wire [46:0] n4480;
  wire [39:0] n4481;
  wire [46:0] n4483;
  wire [3:0] n4485;
  wire n4487;
  wire n4488;
  wire [42:0] n4490;
  wire n4491;
  wire [42:0] n4492;
  wire [42:0] n4493;
  wire [1:0] n4495;
  wire n4497;
  wire n4498;
  wire [40:0] n4500;
  wire n4501;
  wire [40:0] n4502;
  wire [40:0] n4503;
  wire n4505;
  wire n4507;
  wire n4508;
  wire [39:0] n4510;
  wire n4511;
  wire [39:0] n4512;
  wire [39:0] n4513;
  wire [1:0] n4514;
  wire [2:0] n4515;
  wire [3:0] n4516;
  wire [4:0] n4517;
  reg [47:0] n4518;
  reg n4519;
  reg n4520;
  reg [47:0] n4521;
  reg n4522;
  reg n4523;
  reg n4524;
  reg [42:0] n4525;
  reg n4526;
  assign count = scount; //(module output)
  assign r = level0; //(module output)
  /* fplog32.vhdl:2394:16  */
  assign level5_d1 = n4518; // (signal)
  /* fplog32.vhdl:2396:8  */
  assign count4 = n4465; // (signal)
  /* fplog32.vhdl:2396:16  */
  assign count4_d1 = n4519; // (signal)
  /* fplog32.vhdl:2396:27  */
  assign count4_d2 = n4520; // (signal)
  /* fplog32.vhdl:2398:8  */
  assign level4 = n4468; // (signal)
  /* fplog32.vhdl:2398:16  */
  assign level4_d1 = n4521; // (signal)
  /* fplog32.vhdl:2400:8  */
  assign count3 = n4476; // (signal)
  /* fplog32.vhdl:2400:16  */
  assign count3_d1 = n4522; // (signal)
  /* fplog32.vhdl:2400:27  */
  assign count3_d2 = n4523; // (signal)
  /* fplog32.vhdl:2402:8  */
  assign level3 = n4480; // (signal)
  /* fplog32.vhdl:2404:8  */
  assign count2 = n4488; // (signal)
  /* fplog32.vhdl:2404:16  */
  assign count2_d1 = n4524; // (signal)
  /* fplog32.vhdl:2406:8  */
  assign level2 = n4492; // (signal)
  /* fplog32.vhdl:2406:16  */
  assign level2_d1 = n4525; // (signal)
  /* fplog32.vhdl:2408:8  */
  assign count1 = n4498; // (signal)
  /* fplog32.vhdl:2408:16  */
  assign count1_d1 = n4526; // (signal)
  /* fplog32.vhdl:2410:8  */
  assign level1 = n4502; // (signal)
  /* fplog32.vhdl:2412:8  */
  assign count0 = n4508; // (signal)
  /* fplog32.vhdl:2414:8  */
  assign level0 = n4512; // (signal)
  /* fplog32.vhdl:2416:8  */
  assign scount = n4517; // (signal)
  /* fplog32.vhdl:2434:31  */
  assign n4462 = level5_d1[47:32]; // extract
  /* fplog32.vhdl:2434:46  */
  assign n4464 = n4462 == 16'b0000000000000000;
  /* fplog32.vhdl:2434:17  */
  assign n4465 = n4464 ? 1'b1 : 1'b0;
  /* fplog32.vhdl:2435:47  */
  assign n4467 = ~count4;
  /* fplog32.vhdl:2435:36  */
  assign n4468 = n4467 ? level5_d1 : n4471;
  /* fplog32.vhdl:2435:66  */
  assign n4469 = level5_d1[31:0]; // extract
  /* fplog32.vhdl:2435:80  */
  assign n4471 = {n4469, 16'b0000000000000000};
  /* fplog32.vhdl:2437:28  */
  assign n4473 = level4[47:40]; // extract
  /* fplog32.vhdl:2437:43  */
  assign n4475 = n4473 == 8'b00000000;
  /* fplog32.vhdl:2437:17  */
  assign n4476 = n4475 ? 1'b1 : 1'b0;
  /* fplog32.vhdl:2438:22  */
  assign n4478 = level4_d1[47:1]; // extract
  /* fplog32.vhdl:2438:50  */
  assign n4479 = ~count3_d1;
  /* fplog32.vhdl:2438:36  */
  assign n4480 = n4479 ? n4478 : n4483;
  /* fplog32.vhdl:2438:69  */
  assign n4481 = level4_d1[39:0]; // extract
  /* fplog32.vhdl:2438:83  */
  assign n4483 = {n4481, 7'b0000000};
  /* fplog32.vhdl:2440:28  */
  assign n4485 = level3[46:43]; // extract
  /* fplog32.vhdl:2440:43  */
  assign n4487 = n4485 == 4'b0000;
  /* fplog32.vhdl:2440:17  */
  assign n4488 = n4487 ? 1'b1 : 1'b0;
  /* fplog32.vhdl:2441:19  */
  assign n4490 = level3[46:4]; // extract
  /* fplog32.vhdl:2441:44  */
  assign n4491 = ~count2;
  /* fplog32.vhdl:2441:33  */
  assign n4492 = n4491 ? n4490 : n4493;
  /* fplog32.vhdl:2441:60  */
  assign n4493 = level3[42:0]; // extract
  /* fplog32.vhdl:2443:28  */
  assign n4495 = level2[42:41]; // extract
  /* fplog32.vhdl:2443:43  */
  assign n4497 = n4495 == 2'b00;
  /* fplog32.vhdl:2443:17  */
  assign n4498 = n4497 ? 1'b1 : 1'b0;
  /* fplog32.vhdl:2444:22  */
  assign n4500 = level2_d1[42:2]; // extract
  /* fplog32.vhdl:2444:50  */
  assign n4501 = ~count1_d1;
  /* fplog32.vhdl:2444:36  */
  assign n4502 = n4501 ? n4500 : n4503;
  /* fplog32.vhdl:2444:69  */
  assign n4503 = level2_d1[40:0]; // extract
  /* fplog32.vhdl:2446:28  */
  assign n4505 = level1[40]; // extract
  /* fplog32.vhdl:2446:43  */
  assign n4507 = n4505 == 1'b0;
  /* fplog32.vhdl:2446:17  */
  assign n4508 = n4507 ? 1'b1 : 1'b0;
  /* fplog32.vhdl:2447:19  */
  assign n4510 = level1[40:1]; // extract
  /* fplog32.vhdl:2447:44  */
  assign n4511 = ~count0;
  /* fplog32.vhdl:2447:33  */
  assign n4512 = n4511 ? n4510 : n4513;
  /* fplog32.vhdl:2447:60  */
  assign n4513 = level1[39:0]; // extract
  /* fplog32.vhdl:2450:24  */
  assign n4514 = {count4_d2, count3_d2};
  /* fplog32.vhdl:2450:36  */
  assign n4515 = {n4514, count2_d1};
  /* fplog32.vhdl:2450:48  */
  assign n4516 = {n4515, count1_d1};
  /* fplog32.vhdl:2450:60  */
  assign n4517 = {n4516, count0};
  /* fplog32.vhdl:2421:10  */
  always @(posedge clk)
    n4518 <= level5;
  /* fplog32.vhdl:2421:10  */
  always @(posedge clk)
    n4519 <= count4;
  /* fplog32.vhdl:2421:10  */
  always @(posedge clk)
    n4520 <= count4_d1;
  /* fplog32.vhdl:2421:10  */
  always @(posedge clk)
    n4521 <= level4;
  /* fplog32.vhdl:2421:10  */
  always @(posedge clk)
    n4522 <= count3;
  /* fplog32.vhdl:2421:10  */
  always @(posedge clk)
    n4523 <= count3_d1;
  /* fplog32.vhdl:2421:10  */
  always @(posedge clk)
    n4524 <= count2;
  /* fplog32.vhdl:2421:10  */
  always @(posedge clk)
    n4525 <= level2;
  /* fplog32.vhdl:2421:10  */
  always @(posedge clk)
    n4526 <= count1;
endmodule

module intadder_48_freq500_uid43
  (input  clk,
   input  [47:0] x,
   input  [47:0] y,
   input  cin,
   output [47:0] r);
  wire cin_0;
  wire cin_0_d1;
  wire cin_0_d2;
  wire cin_0_d3;
  wire cin_0_d4;
  wire cin_0_d5;
  wire cin_0_d6;
  wire cin_0_d7;
  wire cin_0_d8;
  wire [3:0] x_0;
  wire [3:0] x_0_d1;
  wire [3:0] x_0_d2;
  wire [3:0] x_0_d3;
  wire [3:0] x_0_d4;
  wire [3:0] x_0_d5;
  wire [3:0] x_0_d6;
  wire [3:0] x_0_d7;
  wire [3:0] y_0;
  wire [3:0] y_0_d1;
  wire [3:0] s_0;
  wire [2:0] r_0;
  wire cin_1;
  wire [45:0] x_1;
  wire [45:0] x_1_d1;
  wire [45:0] x_1_d2;
  wire [45:0] x_1_d3;
  wire [45:0] x_1_d4;
  wire [45:0] x_1_d5;
  wire [45:0] x_1_d6;
  wire [45:0] x_1_d7;
  wire [45:0] y_1;
  wire [45:0] y_1_d1;
  wire [45:0] s_1;
  wire [44:0] r_1;
  wire [2:0] n4400;
  wire [3:0] n4402;
  wire [2:0] n4403;
  wire [3:0] n4405;
  wire [3:0] n4406;
  wire [3:0] n4407;
  wire [3:0] n4408;
  wire [2:0] n4409;
  wire n4410;
  wire [44:0] n4411;
  wire [45:0] n4413;
  wire [44:0] n4414;
  wire [45:0] n4416;
  wire [45:0] n4417;
  wire [45:0] n4418;
  wire [45:0] n4419;
  wire [44:0] n4420;
  wire [47:0] n4421;
  reg n4422;
  reg n4423;
  reg n4424;
  reg n4425;
  reg n4426;
  reg n4427;
  reg n4428;
  reg n4429;
  reg [3:0] n4430;
  reg [3:0] n4431;
  reg [3:0] n4432;
  reg [3:0] n4433;
  reg [3:0] n4434;
  reg [3:0] n4435;
  reg [3:0] n4436;
  reg [3:0] n4437;
  reg [45:0] n4438;
  reg [45:0] n4439;
  reg [45:0] n4440;
  reg [45:0] n4441;
  reg [45:0] n4442;
  reg [45:0] n4443;
  reg [45:0] n4444;
  reg [45:0] n4445;
  assign r = n4421; //(module output)
  /* fplog32.vhdl:2300:15  */
  assign cin_0_d1 = n4422; // (signal)
  /* fplog32.vhdl:2300:25  */
  assign cin_0_d2 = n4423; // (signal)
  /* fplog32.vhdl:2300:35  */
  assign cin_0_d3 = n4424; // (signal)
  /* fplog32.vhdl:2300:45  */
  assign cin_0_d4 = n4425; // (signal)
  /* fplog32.vhdl:2300:55  */
  assign cin_0_d5 = n4426; // (signal)
  /* fplog32.vhdl:2300:65  */
  assign cin_0_d6 = n4427; // (signal)
  /* fplog32.vhdl:2300:75  */
  assign cin_0_d7 = n4428; // (signal)
  /* fplog32.vhdl:2300:85  */
  assign cin_0_d8 = n4429; // (signal)
  /* fplog32.vhdl:2302:8  */
  assign x_0 = n4402; // (signal)
  /* fplog32.vhdl:2302:13  */
  assign x_0_d1 = n4430; // (signal)
  /* fplog32.vhdl:2302:21  */
  assign x_0_d2 = n4431; // (signal)
  /* fplog32.vhdl:2302:29  */
  assign x_0_d3 = n4432; // (signal)
  /* fplog32.vhdl:2302:37  */
  assign x_0_d4 = n4433; // (signal)
  /* fplog32.vhdl:2302:45  */
  assign x_0_d5 = n4434; // (signal)
  /* fplog32.vhdl:2302:53  */
  assign x_0_d6 = n4435; // (signal)
  /* fplog32.vhdl:2302:61  */
  assign x_0_d7 = n4436; // (signal)
  /* fplog32.vhdl:2304:8  */
  assign y_0 = n4405; // (signal)
  /* fplog32.vhdl:2304:13  */
  assign y_0_d1 = n4437; // (signal)
  /* fplog32.vhdl:2306:8  */
  assign s_0 = n4408; // (signal)
  /* fplog32.vhdl:2308:8  */
  assign r_0 = n4409; // (signal)
  /* fplog32.vhdl:2310:8  */
  assign cin_1 = n4410; // (signal)
  /* fplog32.vhdl:2312:8  */
  assign x_1 = n4413; // (signal)
  /* fplog32.vhdl:2312:13  */
  assign x_1_d1 = n4438; // (signal)
  /* fplog32.vhdl:2312:21  */
  assign x_1_d2 = n4439; // (signal)
  /* fplog32.vhdl:2312:29  */
  assign x_1_d3 = n4440; // (signal)
  /* fplog32.vhdl:2312:37  */
  assign x_1_d4 = n4441; // (signal)
  /* fplog32.vhdl:2312:45  */
  assign x_1_d5 = n4442; // (signal)
  /* fplog32.vhdl:2312:53  */
  assign x_1_d6 = n4443; // (signal)
  /* fplog32.vhdl:2312:61  */
  assign x_1_d7 = n4444; // (signal)
  /* fplog32.vhdl:2314:8  */
  assign y_1 = n4416; // (signal)
  /* fplog32.vhdl:2314:13  */
  assign y_1_d1 = n4445; // (signal)
  /* fplog32.vhdl:2316:8  */
  assign s_1 = n4419; // (signal)
  /* fplog32.vhdl:2318:8  */
  assign r_1 = n4420; // (signal)
  /* fplog32.vhdl:2351:18  */
  assign n4400 = x[2:0]; // extract
  /* fplog32.vhdl:2351:15  */
  assign n4402 = {1'b0, n4400};
  /* fplog32.vhdl:2352:18  */
  assign n4403 = y[2:0]; // extract
  /* fplog32.vhdl:2352:15  */
  assign n4405 = {1'b0, n4403};
  /* fplog32.vhdl:2353:18  */
  assign n4406 = x_0_d7 + y_0_d1;
  /* fplog32.vhdl:2353:27  */
  assign n4407 = {3'b0, cin_0_d8};  //  uext
  /* fplog32.vhdl:2353:27  */
  assign n4408 = n4406 + n4407;
  /* fplog32.vhdl:2354:14  */
  assign n4409 = s_0[2:0]; // extract
  /* fplog32.vhdl:2355:16  */
  assign n4410 = s_0[3]; // extract
  /* fplog32.vhdl:2356:18  */
  assign n4411 = x[47:3]; // extract
  /* fplog32.vhdl:2356:15  */
  assign n4413 = {1'b0, n4411};
  /* fplog32.vhdl:2357:18  */
  assign n4414 = y[47:3]; // extract
  /* fplog32.vhdl:2357:15  */
  assign n4416 = {1'b0, n4414};
  /* fplog32.vhdl:2358:18  */
  assign n4417 = x_1_d7 + y_1_d1;
  /* fplog32.vhdl:2358:27  */
  assign n4418 = {45'b0, cin_1};  //  uext
  /* fplog32.vhdl:2358:27  */
  assign n4419 = n4417 + n4418;
  /* fplog32.vhdl:2359:14  */
  assign n4420 = s_1[44:0]; // extract
  /* fplog32.vhdl:2360:13  */
  assign n4421 = {r_1, r_0};
  /* fplog32.vhdl:2323:10  */
  always @(posedge clk)
    n4422 <= cin_0;
  /* fplog32.vhdl:2323:10  */
  always @(posedge clk)
    n4423 <= cin_0_d1;
  /* fplog32.vhdl:2323:10  */
  always @(posedge clk)
    n4424 <= cin_0_d2;
  /* fplog32.vhdl:2323:10  */
  always @(posedge clk)
    n4425 <= cin_0_d3;
  /* fplog32.vhdl:2323:10  */
  always @(posedge clk)
    n4426 <= cin_0_d4;
  /* fplog32.vhdl:2323:10  */
  always @(posedge clk)
    n4427 <= cin_0_d5;
  /* fplog32.vhdl:2323:10  */
  always @(posedge clk)
    n4428 <= cin_0_d6;
  /* fplog32.vhdl:2323:10  */
  always @(posedge clk)
    n4429 <= cin_0_d7;
  /* fplog32.vhdl:2323:10  */
  always @(posedge clk)
    n4430 <= x_0;
  /* fplog32.vhdl:2323:10  */
  always @(posedge clk)
    n4431 <= x_0_d1;
  /* fplog32.vhdl:2323:10  */
  always @(posedge clk)
    n4432 <= x_0_d2;
  /* fplog32.vhdl:2323:10  */
  always @(posedge clk)
    n4433 <= x_0_d3;
  /* fplog32.vhdl:2323:10  */
  always @(posedge clk)
    n4434 <= x_0_d4;
  /* fplog32.vhdl:2323:10  */
  always @(posedge clk)
    n4435 <= x_0_d5;
  /* fplog32.vhdl:2323:10  */
  always @(posedge clk)
    n4436 <= x_0_d6;
  /* fplog32.vhdl:2323:10  */
  always @(posedge clk)
    n4437 <= y_0;
  /* fplog32.vhdl:2323:10  */
  always @(posedge clk)
    n4438 <= x_1;
  /* fplog32.vhdl:2323:10  */
  always @(posedge clk)
    n4439 <= x_1_d1;
  /* fplog32.vhdl:2323:10  */
  always @(posedge clk)
    n4440 <= x_1_d2;
  /* fplog32.vhdl:2323:10  */
  always @(posedge clk)
    n4441 <= x_1_d3;
  /* fplog32.vhdl:2323:10  */
  always @(posedge clk)
    n4442 <= x_1_d4;
  /* fplog32.vhdl:2323:10  */
  always @(posedge clk)
    n4443 <= x_1_d5;
  /* fplog32.vhdl:2323:10  */
  always @(posedge clk)
    n4444 <= x_1_d6;
  /* fplog32.vhdl:2323:10  */
  always @(posedge clk)
    n4445 <= y_1;
endmodule

module fixrealkcm_freq500_uid31
  (input  clk,
   input  [7:0] x,
   output [34:0] r);
  wire [4:0] fixrealkcm_freq500_uid31_a0;
  wire [34:0] fixrealkcm_freq500_uid31_t0;
  wire [34:0] fixrealkcm_freq500_uid31_t0_copy35;
  wire [34:0] fixrealkcm_freq500_uid31_t0_copy35_d1;
  wire bh32_w0_0;
  wire bh32_w1_0;
  wire bh32_w2_0;
  wire bh32_w3_0;
  wire bh32_w4_0;
  wire bh32_w5_0;
  wire bh32_w6_0;
  wire bh32_w7_0;
  wire bh32_w8_0;
  wire bh32_w9_0;
  wire bh32_w10_0;
  wire bh32_w11_0;
  wire bh32_w12_0;
  wire bh32_w13_0;
  wire bh32_w14_0;
  wire bh32_w15_0;
  wire bh32_w16_0;
  wire bh32_w17_0;
  wire bh32_w18_0;
  wire bh32_w19_0;
  wire bh32_w20_0;
  wire bh32_w21_0;
  wire bh32_w22_0;
  wire bh32_w23_0;
  wire bh32_w24_0;
  wire bh32_w25_0;
  wire bh32_w26_0;
  wire bh32_w27_0;
  wire bh32_w28_0;
  wire bh32_w29_0;
  wire bh32_w30_0;
  wire bh32_w31_0;
  wire bh32_w32_0;
  wire bh32_w33_0;
  wire bh32_w34_0;
  wire [2:0] fixrealkcm_freq500_uid31_a1;
  wire [29:0] fixrealkcm_freq500_uid31_t1;
  wire [29:0] fixrealkcm_freq500_uid31_t1_copy38;
  wire [29:0] fixrealkcm_freq500_uid31_t1_copy38_d1;
  wire bh32_w0_1;
  wire bh32_w1_1;
  wire bh32_w2_1;
  wire bh32_w3_1;
  wire bh32_w4_1;
  wire bh32_w5_1;
  wire bh32_w6_1;
  wire bh32_w7_1;
  wire bh32_w8_1;
  wire bh32_w9_1;
  wire bh32_w10_1;
  wire bh32_w11_1;
  wire bh32_w12_1;
  wire bh32_w13_1;
  wire bh32_w14_1;
  wire bh32_w15_1;
  wire bh32_w16_1;
  wire bh32_w17_1;
  wire bh32_w18_1;
  wire bh32_w19_1;
  wire bh32_w20_1;
  wire bh32_w21_1;
  wire bh32_w22_1;
  wire bh32_w23_1;
  wire bh32_w24_1;
  wire bh32_w25_1;
  wire bh32_w26_1;
  wire bh32_w27_1;
  wire bh32_w28_1;
  wire bh32_w29_1;
  wire [34:0] bitheapfinaladd_bh32_in0;
  wire [34:0] bitheapfinaladd_bh32_in1;
  wire bitheapfinaladd_bh32_cin;
  wire [34:0] bitheapfinaladd_bh32_out;
  wire [34:0] bitheapresult_bh32;
  wire [34:0] outres;
  wire [4:0] n4226;
  wire [34:0] fixrealkcm_freq500_uid31_table0_n4227;
  wire n4230;
  wire n4231;
  wire n4232;
  wire n4233;
  wire n4234;
  wire n4235;
  wire n4236;
  wire n4237;
  wire n4238;
  wire n4239;
  wire n4240;
  wire n4241;
  wire n4242;
  wire n4243;
  wire n4244;
  wire n4245;
  wire n4246;
  wire n4247;
  wire n4248;
  wire n4249;
  wire n4250;
  wire n4251;
  wire n4252;
  wire n4253;
  wire n4254;
  wire n4255;
  wire n4256;
  wire n4257;
  wire n4258;
  wire n4259;
  wire n4260;
  wire n4261;
  wire n4262;
  wire n4263;
  wire n4264;
  wire [2:0] n4265;
  wire [29:0] fixrealkcm_freq500_uid31_table1_n4266;
  wire n4269;
  wire n4270;
  wire n4271;
  wire n4272;
  wire n4273;
  wire n4274;
  wire n4275;
  wire n4276;
  wire n4277;
  wire n4278;
  wire n4279;
  wire n4280;
  wire n4281;
  wire n4282;
  wire n4283;
  wire n4284;
  wire n4285;
  wire n4286;
  wire n4287;
  wire n4288;
  wire n4289;
  wire n4290;
  wire n4291;
  wire n4292;
  wire n4293;
  wire n4294;
  wire n4295;
  wire n4296;
  wire n4297;
  wire n4298;
  wire [1:0] n4300;
  wire [2:0] n4301;
  wire [3:0] n4302;
  wire [4:0] n4303;
  wire [5:0] n4304;
  wire [6:0] n4305;
  wire [7:0] n4306;
  wire [8:0] n4307;
  wire [9:0] n4308;
  wire [10:0] n4309;
  wire [11:0] n4310;
  wire [12:0] n4311;
  wire [13:0] n4312;
  wire [14:0] n4313;
  wire [15:0] n4314;
  wire [16:0] n4315;
  wire [17:0] n4316;
  wire [18:0] n4317;
  wire [19:0] n4318;
  wire [20:0] n4319;
  wire [21:0] n4320;
  wire [22:0] n4321;
  wire [23:0] n4322;
  wire [24:0] n4323;
  wire [25:0] n4324;
  wire [26:0] n4325;
  wire [27:0] n4326;
  wire [28:0] n4327;
  wire [29:0] n4328;
  wire [30:0] n4329;
  wire [31:0] n4330;
  wire [32:0] n4331;
  wire [33:0] n4332;
  wire [34:0] n4333;
  wire [5:0] n4335;
  wire [6:0] n4336;
  wire [7:0] n4337;
  wire [8:0] n4338;
  wire [9:0] n4339;
  wire [10:0] n4340;
  wire [11:0] n4341;
  wire [12:0] n4342;
  wire [13:0] n4343;
  wire [14:0] n4344;
  wire [15:0] n4345;
  wire [16:0] n4346;
  wire [17:0] n4347;
  wire [18:0] n4348;
  wire [19:0] n4349;
  wire [20:0] n4350;
  wire [21:0] n4351;
  wire [22:0] n4352;
  wire [23:0] n4353;
  wire [24:0] n4354;
  wire [25:0] n4355;
  wire [26:0] n4356;
  wire [27:0] n4357;
  wire [28:0] n4358;
  wire [29:0] n4359;
  wire [30:0] n4360;
  wire [31:0] n4361;
  wire [32:0] n4362;
  wire [33:0] n4363;
  wire [34:0] n4364;
  wire [34:0] bitheapfinaladd_bh32_n4366;
  reg [34:0] n4369;
  reg [29:0] n4370;
  assign r = outres; //(module output)
  /* fplog32.vhdl:2010:8  */
  assign fixrealkcm_freq500_uid31_a0 = n4226; // (signal)
  /* fplog32.vhdl:2012:8  */
  assign fixrealkcm_freq500_uid31_t0 = fixrealkcm_freq500_uid31_t0_copy35_d1; // (signal)
  /* fplog32.vhdl:2014:8  */
  assign fixrealkcm_freq500_uid31_t0_copy35 = fixrealkcm_freq500_uid31_table0_n4227; // (signal)
  /* fplog32.vhdl:2014:44  */
  assign fixrealkcm_freq500_uid31_t0_copy35_d1 = n4369; // (signal)
  /* fplog32.vhdl:2016:8  */
  assign bh32_w0_0 = n4230; // (signal)
  /* fplog32.vhdl:2018:8  */
  assign bh32_w1_0 = n4231; // (signal)
  /* fplog32.vhdl:2020:8  */
  assign bh32_w2_0 = n4232; // (signal)
  /* fplog32.vhdl:2022:8  */
  assign bh32_w3_0 = n4233; // (signal)
  /* fplog32.vhdl:2024:8  */
  assign bh32_w4_0 = n4234; // (signal)
  /* fplog32.vhdl:2026:8  */
  assign bh32_w5_0 = n4235; // (signal)
  /* fplog32.vhdl:2028:8  */
  assign bh32_w6_0 = n4236; // (signal)
  /* fplog32.vhdl:2030:8  */
  assign bh32_w7_0 = n4237; // (signal)
  /* fplog32.vhdl:2032:8  */
  assign bh32_w8_0 = n4238; // (signal)
  /* fplog32.vhdl:2034:8  */
  assign bh32_w9_0 = n4239; // (signal)
  /* fplog32.vhdl:2036:8  */
  assign bh32_w10_0 = n4240; // (signal)
  /* fplog32.vhdl:2038:8  */
  assign bh32_w11_0 = n4241; // (signal)
  /* fplog32.vhdl:2040:8  */
  assign bh32_w12_0 = n4242; // (signal)
  /* fplog32.vhdl:2042:8  */
  assign bh32_w13_0 = n4243; // (signal)
  /* fplog32.vhdl:2044:8  */
  assign bh32_w14_0 = n4244; // (signal)
  /* fplog32.vhdl:2046:8  */
  assign bh32_w15_0 = n4245; // (signal)
  /* fplog32.vhdl:2048:8  */
  assign bh32_w16_0 = n4246; // (signal)
  /* fplog32.vhdl:2050:8  */
  assign bh32_w17_0 = n4247; // (signal)
  /* fplog32.vhdl:2052:8  */
  assign bh32_w18_0 = n4248; // (signal)
  /* fplog32.vhdl:2054:8  */
  assign bh32_w19_0 = n4249; // (signal)
  /* fplog32.vhdl:2056:8  */
  assign bh32_w20_0 = n4250; // (signal)
  /* fplog32.vhdl:2058:8  */
  assign bh32_w21_0 = n4251; // (signal)
  /* fplog32.vhdl:2060:8  */
  assign bh32_w22_0 = n4252; // (signal)
  /* fplog32.vhdl:2062:8  */
  assign bh32_w23_0 = n4253; // (signal)
  /* fplog32.vhdl:2064:8  */
  assign bh32_w24_0 = n4254; // (signal)
  /* fplog32.vhdl:2066:8  */
  assign bh32_w25_0 = n4255; // (signal)
  /* fplog32.vhdl:2068:8  */
  assign bh32_w26_0 = n4256; // (signal)
  /* fplog32.vhdl:2070:8  */
  assign bh32_w27_0 = n4257; // (signal)
  /* fplog32.vhdl:2072:8  */
  assign bh32_w28_0 = n4258; // (signal)
  /* fplog32.vhdl:2074:8  */
  assign bh32_w29_0 = n4259; // (signal)
  /* fplog32.vhdl:2076:8  */
  assign bh32_w30_0 = n4260; // (signal)
  /* fplog32.vhdl:2078:8  */
  assign bh32_w31_0 = n4261; // (signal)
  /* fplog32.vhdl:2080:8  */
  assign bh32_w32_0 = n4262; // (signal)
  /* fplog32.vhdl:2082:8  */
  assign bh32_w33_0 = n4263; // (signal)
  /* fplog32.vhdl:2253:35  */
  assign bh32_w34_0 = n4264; // (signal)
  /* fplog32.vhdl:2086:8  */
  assign fixrealkcm_freq500_uid31_a1 = n4265; // (signal)
  /* fplog32.vhdl:2088:8  */
  assign fixrealkcm_freq500_uid31_t1 = fixrealkcm_freq500_uid31_t1_copy38_d1; // (signal)
  /* fplog32.vhdl:2090:8  */
  assign fixrealkcm_freq500_uid31_t1_copy38 = fixrealkcm_freq500_uid31_table1_n4266; // (signal)
  /* fplog32.vhdl:2090:44  */
  assign fixrealkcm_freq500_uid31_t1_copy38_d1 = n4370; // (signal)
  /* fplog32.vhdl:2092:8  */
  assign bh32_w0_1 = n4269; // (signal)
  /* fplog32.vhdl:2094:8  */
  assign bh32_w1_1 = n4270; // (signal)
  /* fplog32.vhdl:2096:8  */
  assign bh32_w2_1 = n4271; // (signal)
  /* fplog32.vhdl:2098:8  */
  assign bh32_w3_1 = n4272; // (signal)
  /* fplog32.vhdl:2100:8  */
  assign bh32_w4_1 = n4273; // (signal)
  /* fplog32.vhdl:2102:8  */
  assign bh32_w5_1 = n4274; // (signal)
  /* fplog32.vhdl:2104:8  */
  assign bh32_w6_1 = n4275; // (signal)
  /* fplog32.vhdl:2106:8  */
  assign bh32_w7_1 = n4276; // (signal)
  /* fplog32.vhdl:2108:8  */
  assign bh32_w8_1 = n4277; // (signal)
  /* fplog32.vhdl:2110:8  */
  assign bh32_w9_1 = n4278; // (signal)
  /* fplog32.vhdl:2112:8  */
  assign bh32_w10_1 = n4279; // (signal)
  /* fplog32.vhdl:2114:8  */
  assign bh32_w11_1 = n4280; // (signal)
  /* fplog32.vhdl:2116:8  */
  assign bh32_w12_1 = n4281; // (signal)
  /* fplog32.vhdl:2118:8  */
  assign bh32_w13_1 = n4282; // (signal)
  /* fplog32.vhdl:2120:8  */
  assign bh32_w14_1 = n4283; // (signal)
  /* fplog32.vhdl:2122:8  */
  assign bh32_w15_1 = n4284; // (signal)
  /* fplog32.vhdl:2124:8  */
  assign bh32_w16_1 = n4285; // (signal)
  /* fplog32.vhdl:2126:8  */
  assign bh32_w17_1 = n4286; // (signal)
  /* fplog32.vhdl:2128:8  */
  assign bh32_w18_1 = n4287; // (signal)
  /* fplog32.vhdl:2130:8  */
  assign bh32_w19_1 = n4288; // (signal)
  /* fplog32.vhdl:2132:8  */
  assign bh32_w20_1 = n4289; // (signal)
  /* fplog32.vhdl:2134:8  */
  assign bh32_w21_1 = n4290; // (signal)
  /* fplog32.vhdl:2136:8  */
  assign bh32_w22_1 = n4291; // (signal)
  /* fplog32.vhdl:2138:8  */
  assign bh32_w23_1 = n4292; // (signal)
  /* fplog32.vhdl:2140:8  */
  assign bh32_w24_1 = n4293; // (signal)
  /* fplog32.vhdl:2142:8  */
  assign bh32_w25_1 = n4294; // (signal)
  /* fplog32.vhdl:2144:8  */
  assign bh32_w26_1 = n4295; // (signal)
  /* fplog32.vhdl:2146:8  */
  assign bh32_w27_1 = n4296; // (signal)
  /* fplog32.vhdl:2148:8  */
  assign bh32_w28_1 = n4297; // (signal)
  /* fplog32.vhdl:2150:8  */
  assign bh32_w29_1 = n4298; // (signal)
  /* fplog32.vhdl:2152:8  */
  assign bitheapfinaladd_bh32_in0 = n4333; // (signal)
  /* fplog32.vhdl:2154:8  */
  assign bitheapfinaladd_bh32_in1 = n4364; // (signal)
  /* fplog32.vhdl:2156:8  */
  assign bitheapfinaladd_bh32_cin = 1'b0; // (signal)
  /* fplog32.vhdl:2158:8  */
  assign bitheapfinaladd_bh32_out = bitheapfinaladd_bh32_n4366; // (signal)
  /* fplog32.vhdl:2160:8  */
  assign bitheapresult_bh32 = bitheapfinaladd_bh32_out; // (signal)
  /* fplog32.vhdl:2162:8  */
  assign outres = bitheapresult_bh32; // (signal)
  /* fplog32.vhdl:2173:36  */
  assign n4226 = x[7:3]; // extract
  /* fplog32.vhdl:2174:4  */
  fixrealkcm_freq500_uid31_t0_freq500_uid34 fixrealkcm_freq500_uid31_table0 (
    .x(fixrealkcm_freq500_uid31_a0),
    .y(fixrealkcm_freq500_uid31_table0_n4227));
  /* fplog32.vhdl:2178:44  */
  assign n4230 = fixrealkcm_freq500_uid31_t0[0]; // extract
  /* fplog32.vhdl:2179:44  */
  assign n4231 = fixrealkcm_freq500_uid31_t0[1]; // extract
  /* fplog32.vhdl:2180:44  */
  assign n4232 = fixrealkcm_freq500_uid31_t0[2]; // extract
  /* fplog32.vhdl:2181:44  */
  assign n4233 = fixrealkcm_freq500_uid31_t0[3]; // extract
  /* fplog32.vhdl:2182:44  */
  assign n4234 = fixrealkcm_freq500_uid31_t0[4]; // extract
  /* fplog32.vhdl:2183:44  */
  assign n4235 = fixrealkcm_freq500_uid31_t0[5]; // extract
  /* fplog32.vhdl:2184:44  */
  assign n4236 = fixrealkcm_freq500_uid31_t0[6]; // extract
  /* fplog32.vhdl:2185:44  */
  assign n4237 = fixrealkcm_freq500_uid31_t0[7]; // extract
  /* fplog32.vhdl:2186:44  */
  assign n4238 = fixrealkcm_freq500_uid31_t0[8]; // extract
  /* fplog32.vhdl:2187:44  */
  assign n4239 = fixrealkcm_freq500_uid31_t0[9]; // extract
  /* fplog32.vhdl:2188:45  */
  assign n4240 = fixrealkcm_freq500_uid31_t0[10]; // extract
  /* fplog32.vhdl:2189:45  */
  assign n4241 = fixrealkcm_freq500_uid31_t0[11]; // extract
  /* fplog32.vhdl:2190:45  */
  assign n4242 = fixrealkcm_freq500_uid31_t0[12]; // extract
  /* fplog32.vhdl:2191:45  */
  assign n4243 = fixrealkcm_freq500_uid31_t0[13]; // extract
  /* fplog32.vhdl:2192:45  */
  assign n4244 = fixrealkcm_freq500_uid31_t0[14]; // extract
  /* fplog32.vhdl:2193:45  */
  assign n4245 = fixrealkcm_freq500_uid31_t0[15]; // extract
  /* fplog32.vhdl:2194:45  */
  assign n4246 = fixrealkcm_freq500_uid31_t0[16]; // extract
  /* fplog32.vhdl:2195:45  */
  assign n4247 = fixrealkcm_freq500_uid31_t0[17]; // extract
  /* fplog32.vhdl:2196:45  */
  assign n4248 = fixrealkcm_freq500_uid31_t0[18]; // extract
  /* fplog32.vhdl:2197:45  */
  assign n4249 = fixrealkcm_freq500_uid31_t0[19]; // extract
  /* fplog32.vhdl:2198:45  */
  assign n4250 = fixrealkcm_freq500_uid31_t0[20]; // extract
  /* fplog32.vhdl:2199:45  */
  assign n4251 = fixrealkcm_freq500_uid31_t0[21]; // extract
  /* fplog32.vhdl:2200:45  */
  assign n4252 = fixrealkcm_freq500_uid31_t0[22]; // extract
  /* fplog32.vhdl:2201:45  */
  assign n4253 = fixrealkcm_freq500_uid31_t0[23]; // extract
  /* fplog32.vhdl:2202:45  */
  assign n4254 = fixrealkcm_freq500_uid31_t0[24]; // extract
  /* fplog32.vhdl:2203:45  */
  assign n4255 = fixrealkcm_freq500_uid31_t0[25]; // extract
  /* fplog32.vhdl:2204:45  */
  assign n4256 = fixrealkcm_freq500_uid31_t0[26]; // extract
  /* fplog32.vhdl:2205:45  */
  assign n4257 = fixrealkcm_freq500_uid31_t0[27]; // extract
  /* fplog32.vhdl:2206:45  */
  assign n4258 = fixrealkcm_freq500_uid31_t0[28]; // extract
  /* fplog32.vhdl:2207:45  */
  assign n4259 = fixrealkcm_freq500_uid31_t0[29]; // extract
  /* fplog32.vhdl:2208:45  */
  assign n4260 = fixrealkcm_freq500_uid31_t0[30]; // extract
  /* fplog32.vhdl:2209:45  */
  assign n4261 = fixrealkcm_freq500_uid31_t0[31]; // extract
  /* fplog32.vhdl:2210:45  */
  assign n4262 = fixrealkcm_freq500_uid31_t0[32]; // extract
  /* fplog32.vhdl:2211:45  */
  assign n4263 = fixrealkcm_freq500_uid31_t0[33]; // extract
  /* fplog32.vhdl:2212:45  */
  assign n4264 = fixrealkcm_freq500_uid31_t0[34]; // extract
  /* fplog32.vhdl:2213:36  */
  assign n4265 = x[2:0]; // extract
  /* fplog32.vhdl:2214:4  */
  fixrealkcm_freq500_uid31_t1_freq500_uid37 fixrealkcm_freq500_uid31_table1 (
    .x(fixrealkcm_freq500_uid31_a1),
    .y(fixrealkcm_freq500_uid31_table1_n4266));
  /* fplog32.vhdl:2218:44  */
  assign n4269 = fixrealkcm_freq500_uid31_t1[0]; // extract
  /* fplog32.vhdl:2219:44  */
  assign n4270 = fixrealkcm_freq500_uid31_t1[1]; // extract
  /* fplog32.vhdl:2220:44  */
  assign n4271 = fixrealkcm_freq500_uid31_t1[2]; // extract
  /* fplog32.vhdl:2221:44  */
  assign n4272 = fixrealkcm_freq500_uid31_t1[3]; // extract
  /* fplog32.vhdl:2222:44  */
  assign n4273 = fixrealkcm_freq500_uid31_t1[4]; // extract
  /* fplog32.vhdl:2223:44  */
  assign n4274 = fixrealkcm_freq500_uid31_t1[5]; // extract
  /* fplog32.vhdl:2224:44  */
  assign n4275 = fixrealkcm_freq500_uid31_t1[6]; // extract
  /* fplog32.vhdl:2225:44  */
  assign n4276 = fixrealkcm_freq500_uid31_t1[7]; // extract
  /* fplog32.vhdl:2226:44  */
  assign n4277 = fixrealkcm_freq500_uid31_t1[8]; // extract
  /* fplog32.vhdl:2227:44  */
  assign n4278 = fixrealkcm_freq500_uid31_t1[9]; // extract
  /* fplog32.vhdl:2228:45  */
  assign n4279 = fixrealkcm_freq500_uid31_t1[10]; // extract
  /* fplog32.vhdl:2229:45  */
  assign n4280 = fixrealkcm_freq500_uid31_t1[11]; // extract
  /* fplog32.vhdl:2230:45  */
  assign n4281 = fixrealkcm_freq500_uid31_t1[12]; // extract
  /* fplog32.vhdl:2231:45  */
  assign n4282 = fixrealkcm_freq500_uid31_t1[13]; // extract
  /* fplog32.vhdl:2232:45  */
  assign n4283 = fixrealkcm_freq500_uid31_t1[14]; // extract
  /* fplog32.vhdl:2233:45  */
  assign n4284 = fixrealkcm_freq500_uid31_t1[15]; // extract
  /* fplog32.vhdl:2234:45  */
  assign n4285 = fixrealkcm_freq500_uid31_t1[16]; // extract
  /* fplog32.vhdl:2235:45  */
  assign n4286 = fixrealkcm_freq500_uid31_t1[17]; // extract
  /* fplog32.vhdl:2236:45  */
  assign n4287 = fixrealkcm_freq500_uid31_t1[18]; // extract
  /* fplog32.vhdl:2237:45  */
  assign n4288 = fixrealkcm_freq500_uid31_t1[19]; // extract
  /* fplog32.vhdl:2238:45  */
  assign n4289 = fixrealkcm_freq500_uid31_t1[20]; // extract
  /* fplog32.vhdl:2239:45  */
  assign n4290 = fixrealkcm_freq500_uid31_t1[21]; // extract
  /* fplog32.vhdl:2240:45  */
  assign n4291 = fixrealkcm_freq500_uid31_t1[22]; // extract
  /* fplog32.vhdl:2241:45  */
  assign n4292 = fixrealkcm_freq500_uid31_t1[23]; // extract
  /* fplog32.vhdl:2242:45  */
  assign n4293 = fixrealkcm_freq500_uid31_t1[24]; // extract
  /* fplog32.vhdl:2243:45  */
  assign n4294 = fixrealkcm_freq500_uid31_t1[25]; // extract
  /* fplog32.vhdl:2244:45  */
  assign n4295 = fixrealkcm_freq500_uid31_t1[26]; // extract
  /* fplog32.vhdl:2245:45  */
  assign n4296 = fixrealkcm_freq500_uid31_t1[27]; // extract
  /* fplog32.vhdl:2246:45  */
  assign n4297 = fixrealkcm_freq500_uid31_t1[28]; // extract
  /* fplog32.vhdl:2247:45  */
  assign n4298 = fixrealkcm_freq500_uid31_t1[29]; // extract
  /* fplog32.vhdl:2253:48  */
  assign n4300 = {bh32_w34_0, bh32_w33_0};
  /* fplog32.vhdl:2253:61  */
  assign n4301 = {n4300, bh32_w32_0};
  /* fplog32.vhdl:2253:74  */
  assign n4302 = {n4301, bh32_w31_0};
  /* fplog32.vhdl:2253:87  */
  assign n4303 = {n4302, bh32_w30_0};
  /* fplog32.vhdl:2253:100  */
  assign n4304 = {n4303, bh32_w29_1};
  /* fplog32.vhdl:2253:113  */
  assign n4305 = {n4304, bh32_w28_1};
  /* fplog32.vhdl:2253:126  */
  assign n4306 = {n4305, bh32_w27_1};
  /* fplog32.vhdl:2253:139  */
  assign n4307 = {n4306, bh32_w26_1};
  /* fplog32.vhdl:2253:152  */
  assign n4308 = {n4307, bh32_w25_1};
  /* fplog32.vhdl:2253:165  */
  assign n4309 = {n4308, bh32_w24_1};
  /* fplog32.vhdl:2253:178  */
  assign n4310 = {n4309, bh32_w23_1};
  /* fplog32.vhdl:2253:191  */
  assign n4311 = {n4310, bh32_w22_1};
  /* fplog32.vhdl:2253:204  */
  assign n4312 = {n4311, bh32_w21_1};
  /* fplog32.vhdl:2253:217  */
  assign n4313 = {n4312, bh32_w20_1};
  /* fplog32.vhdl:2253:230  */
  assign n4314 = {n4313, bh32_w19_1};
  /* fplog32.vhdl:2253:243  */
  assign n4315 = {n4314, bh32_w18_1};
  /* fplog32.vhdl:2253:256  */
  assign n4316 = {n4315, bh32_w17_1};
  /* fplog32.vhdl:2253:269  */
  assign n4317 = {n4316, bh32_w16_1};
  /* fplog32.vhdl:2253:282  */
  assign n4318 = {n4317, bh32_w15_1};
  /* fplog32.vhdl:2253:295  */
  assign n4319 = {n4318, bh32_w14_1};
  /* fplog32.vhdl:2253:308  */
  assign n4320 = {n4319, bh32_w13_1};
  /* fplog32.vhdl:2253:321  */
  assign n4321 = {n4320, bh32_w12_1};
  /* fplog32.vhdl:2253:334  */
  assign n4322 = {n4321, bh32_w11_1};
  /* fplog32.vhdl:2253:347  */
  assign n4323 = {n4322, bh32_w10_1};
  /* fplog32.vhdl:2253:360  */
  assign n4324 = {n4323, bh32_w9_1};
  /* fplog32.vhdl:2253:372  */
  assign n4325 = {n4324, bh32_w8_1};
  /* fplog32.vhdl:2253:384  */
  assign n4326 = {n4325, bh32_w7_1};
  /* fplog32.vhdl:2253:396  */
  assign n4327 = {n4326, bh32_w6_1};
  /* fplog32.vhdl:2253:408  */
  assign n4328 = {n4327, bh32_w5_1};
  /* fplog32.vhdl:2253:420  */
  assign n4329 = {n4328, bh32_w4_1};
  /* fplog32.vhdl:2253:432  */
  assign n4330 = {n4329, bh32_w3_1};
  /* fplog32.vhdl:2253:444  */
  assign n4331 = {n4330, bh32_w2_1};
  /* fplog32.vhdl:2253:456  */
  assign n4332 = {n4331, bh32_w1_1};
  /* fplog32.vhdl:2253:468  */
  assign n4333 = {n4332, bh32_w0_1};
  /* fplog32.vhdl:2254:60  */
  assign n4335 = {5'b00000, bh32_w29_0};
  /* fplog32.vhdl:2254:73  */
  assign n4336 = {n4335, bh32_w28_0};
  /* fplog32.vhdl:2254:86  */
  assign n4337 = {n4336, bh32_w27_0};
  /* fplog32.vhdl:2254:99  */
  assign n4338 = {n4337, bh32_w26_0};
  /* fplog32.vhdl:2254:112  */
  assign n4339 = {n4338, bh32_w25_0};
  /* fplog32.vhdl:2254:125  */
  assign n4340 = {n4339, bh32_w24_0};
  /* fplog32.vhdl:2254:138  */
  assign n4341 = {n4340, bh32_w23_0};
  /* fplog32.vhdl:2254:151  */
  assign n4342 = {n4341, bh32_w22_0};
  /* fplog32.vhdl:2254:164  */
  assign n4343 = {n4342, bh32_w21_0};
  /* fplog32.vhdl:2254:177  */
  assign n4344 = {n4343, bh32_w20_0};
  /* fplog32.vhdl:2254:190  */
  assign n4345 = {n4344, bh32_w19_0};
  /* fplog32.vhdl:2254:203  */
  assign n4346 = {n4345, bh32_w18_0};
  /* fplog32.vhdl:2254:216  */
  assign n4347 = {n4346, bh32_w17_0};
  /* fplog32.vhdl:2254:229  */
  assign n4348 = {n4347, bh32_w16_0};
  /* fplog32.vhdl:2254:242  */
  assign n4349 = {n4348, bh32_w15_0};
  /* fplog32.vhdl:2254:255  */
  assign n4350 = {n4349, bh32_w14_0};
  /* fplog32.vhdl:2254:268  */
  assign n4351 = {n4350, bh32_w13_0};
  /* fplog32.vhdl:2254:281  */
  assign n4352 = {n4351, bh32_w12_0};
  /* fplog32.vhdl:2254:294  */
  assign n4353 = {n4352, bh32_w11_0};
  /* fplog32.vhdl:2254:307  */
  assign n4354 = {n4353, bh32_w10_0};
  /* fplog32.vhdl:2254:320  */
  assign n4355 = {n4354, bh32_w9_0};
  /* fplog32.vhdl:2254:332  */
  assign n4356 = {n4355, bh32_w8_0};
  /* fplog32.vhdl:2254:344  */
  assign n4357 = {n4356, bh32_w7_0};
  /* fplog32.vhdl:2254:356  */
  assign n4358 = {n4357, bh32_w6_0};
  /* fplog32.vhdl:2254:368  */
  assign n4359 = {n4358, bh32_w5_0};
  /* fplog32.vhdl:2254:380  */
  assign n4360 = {n4359, bh32_w4_0};
  /* fplog32.vhdl:2254:392  */
  assign n4361 = {n4360, bh32_w3_0};
  /* fplog32.vhdl:2254:404  */
  assign n4362 = {n4361, bh32_w2_0};
  /* fplog32.vhdl:2254:416  */
  assign n4363 = {n4362, bh32_w1_0};
  /* fplog32.vhdl:2254:428  */
  assign n4364 = {n4363, bh32_w0_0};
  /* fplog32.vhdl:2257:4  */
  intadder_35_freq500_uid41 bitheapfinaladd_bh32 (
    .clk(clk),
    .x(bitheapfinaladd_bh32_in0),
    .y(bitheapfinaladd_bh32_in1),
    .cin(bitheapfinaladd_bh32_cin),
    .r(bitheapfinaladd_bh32_n4366));
  /* fplog32.vhdl:2167:10  */
  always @(posedge clk)
    n4369 <= fixrealkcm_freq500_uid31_t0_copy35;
  /* fplog32.vhdl:2167:10  */
  always @(posedge clk)
    n4370 <= fixrealkcm_freq500_uid31_t1_copy38;
endmodule

module intadder_40_freq500_uid29
  (input  clk,
   input  [39:0] x,
   input  [39:0] y,
   input  cin,
   output [39:0] r);
  wire cin_1;
  wire cin_1_d1;
  wire cin_1_d2;
  wire cin_1_d3;
  wire cin_1_d4;
  wire cin_1_d5;
  wire cin_1_d6;
  wire cin_1_d7;
  wire [40:0] x_1;
  wire [40:0] x_1_d1;
  wire [40:0] x_1_d2;
  wire [40:0] x_1_d3;
  wire [40:0] x_1_d4;
  wire [40:0] y_1;
  wire [40:0] y_1_d1;
  wire [40:0] s_1;
  wire [39:0] r_1;
  wire [40:0] n4200;
  wire [40:0] n4202;
  wire [40:0] n4203;
  wire [40:0] n4204;
  wire [40:0] n4205;
  wire [39:0] n4206;
  reg n4207;
  reg n4208;
  reg n4209;
  reg n4210;
  reg n4211;
  reg n4212;
  reg n4213;
  reg [40:0] n4214;
  reg [40:0] n4215;
  reg [40:0] n4216;
  reg [40:0] n4217;
  reg [40:0] n4218;
  assign r = r_1; //(module output)
  /* fplog32.vhdl:1879:15  */
  assign cin_1_d1 = n4207; // (signal)
  /* fplog32.vhdl:1879:25  */
  assign cin_1_d2 = n4208; // (signal)
  /* fplog32.vhdl:1879:35  */
  assign cin_1_d3 = n4209; // (signal)
  /* fplog32.vhdl:1879:45  */
  assign cin_1_d4 = n4210; // (signal)
  /* fplog32.vhdl:1879:55  */
  assign cin_1_d5 = n4211; // (signal)
  /* fplog32.vhdl:1879:65  */
  assign cin_1_d6 = n4212; // (signal)
  /* fplog32.vhdl:1879:75  */
  assign cin_1_d7 = n4213; // (signal)
  /* fplog32.vhdl:1881:8  */
  assign x_1 = n4200; // (signal)
  /* fplog32.vhdl:1881:13  */
  assign x_1_d1 = n4214; // (signal)
  /* fplog32.vhdl:1881:21  */
  assign x_1_d2 = n4215; // (signal)
  /* fplog32.vhdl:1881:29  */
  assign x_1_d3 = n4216; // (signal)
  /* fplog32.vhdl:1881:37  */
  assign x_1_d4 = n4217; // (signal)
  /* fplog32.vhdl:1883:8  */
  assign y_1 = n4202; // (signal)
  /* fplog32.vhdl:1883:13  */
  assign y_1_d1 = n4218; // (signal)
  /* fplog32.vhdl:1885:8  */
  assign s_1 = n4205; // (signal)
  /* fplog32.vhdl:1887:8  */
  assign r_1 = n4206; // (signal)
  /* fplog32.vhdl:1908:15  */
  assign n4200 = {1'b0, x};
  /* fplog32.vhdl:1909:15  */
  assign n4202 = {1'b0, y};
  /* fplog32.vhdl:1910:18  */
  assign n4203 = x_1_d4 + y_1_d1;
  /* fplog32.vhdl:1910:27  */
  assign n4204 = {40'b0, cin_1_d7};  //  uext
  /* fplog32.vhdl:1910:27  */
  assign n4205 = n4203 + n4204;
  /* fplog32.vhdl:1911:14  */
  assign n4206 = s_1[39:0]; // extract
  /* fplog32.vhdl:1892:10  */
  always @(posedge clk)
    n4207 <= cin_1;
  /* fplog32.vhdl:1892:10  */
  always @(posedge clk)
    n4208 <= cin_1_d1;
  /* fplog32.vhdl:1892:10  */
  always @(posedge clk)
    n4209 <= cin_1_d2;
  /* fplog32.vhdl:1892:10  */
  always @(posedge clk)
    n4210 <= cin_1_d3;
  /* fplog32.vhdl:1892:10  */
  always @(posedge clk)
    n4211 <= cin_1_d4;
  /* fplog32.vhdl:1892:10  */
  always @(posedge clk)
    n4212 <= cin_1_d5;
  /* fplog32.vhdl:1892:10  */
  always @(posedge clk)
    n4213 <= cin_1_d6;
  /* fplog32.vhdl:1892:10  */
  always @(posedge clk)
    n4214 <= x_1;
  /* fplog32.vhdl:1892:10  */
  always @(posedge clk)
    n4215 <= x_1_d1;
  /* fplog32.vhdl:1892:10  */
  always @(posedge clk)
    n4216 <= x_1_d2;
  /* fplog32.vhdl:1892:10  */
  always @(posedge clk)
    n4217 <= x_1_d3;
  /* fplog32.vhdl:1892:10  */
  always @(posedge clk)
    n4218 <= y_1;
endmodule

module intadder_40_freq500_uid26
  (input  clk,
   input  [39:0] x,
   input  [39:0] y,
   input  cin,
   output [39:0] r);
  wire cin_0;
  wire cin_0_d1;
  wire cin_0_d2;
  wire cin_0_d3;
  wire [39:0] x_0;
  wire [39:0] x_0_d1;
  wire [39:0] y_0;
  wire [39:0] y_0_d1;
  wire [39:0] y_0_d2;
  wire [39:0] s_0;
  wire [38:0] r_0;
  wire cin_1;
  wire [1:0] x_1;
  wire [1:0] x_1_d1;
  wire [1:0] y_1;
  wire [1:0] y_1_d1;
  wire [1:0] y_1_d2;
  wire [1:0] s_1;
  wire r_1;
  wire [38:0] n4151;
  wire [39:0] n4153;
  wire [38:0] n4154;
  wire [39:0] n4156;
  wire [39:0] n4157;
  wire [39:0] n4158;
  wire [39:0] n4159;
  wire [38:0] n4160;
  wire n4161;
  wire n4162;
  wire [1:0] n4164;
  wire n4165;
  wire [1:0] n4167;
  wire [1:0] n4168;
  wire [1:0] n4169;
  wire [1:0] n4170;
  wire n4171;
  wire [39:0] n4172;
  reg n4173;
  reg n4174;
  reg n4175;
  reg [39:0] n4176;
  reg [39:0] n4177;
  reg [39:0] n4178;
  reg [1:0] n4179;
  reg [1:0] n4180;
  reg [1:0] n4181;
  assign r = n4172; //(module output)
  /* fplog32.vhdl:1799:15  */
  assign cin_0_d1 = n4173; // (signal)
  /* fplog32.vhdl:1799:25  */
  assign cin_0_d2 = n4174; // (signal)
  /* fplog32.vhdl:1799:35  */
  assign cin_0_d3 = n4175; // (signal)
  /* fplog32.vhdl:1801:8  */
  assign x_0 = n4153; // (signal)
  /* fplog32.vhdl:1801:13  */
  assign x_0_d1 = n4176; // (signal)
  /* fplog32.vhdl:1803:8  */
  assign y_0 = n4156; // (signal)
  /* fplog32.vhdl:1803:13  */
  assign y_0_d1 = n4177; // (signal)
  /* fplog32.vhdl:1803:21  */
  assign y_0_d2 = n4178; // (signal)
  /* fplog32.vhdl:1805:8  */
  assign s_0 = n4159; // (signal)
  /* fplog32.vhdl:1807:8  */
  assign r_0 = n4160; // (signal)
  /* fplog32.vhdl:1809:8  */
  assign cin_1 = n4161; // (signal)
  /* fplog32.vhdl:1811:8  */
  assign x_1 = n4164; // (signal)
  /* fplog32.vhdl:1811:13  */
  assign x_1_d1 = n4179; // (signal)
  /* fplog32.vhdl:1813:8  */
  assign y_1 = n4167; // (signal)
  /* fplog32.vhdl:1813:13  */
  assign y_1_d1 = n4180; // (signal)
  /* fplog32.vhdl:1813:21  */
  assign y_1_d2 = n4181; // (signal)
  /* fplog32.vhdl:1815:8  */
  assign s_1 = n4170; // (signal)
  /* fplog32.vhdl:1817:8  */
  assign r_1 = n4171; // (signal)
  /* fplog32.vhdl:1835:18  */
  assign n4151 = x[38:0]; // extract
  /* fplog32.vhdl:1835:15  */
  assign n4153 = {1'b0, n4151};
  /* fplog32.vhdl:1836:18  */
  assign n4154 = y[38:0]; // extract
  /* fplog32.vhdl:1836:15  */
  assign n4156 = {1'b0, n4154};
  /* fplog32.vhdl:1837:18  */
  assign n4157 = x_0_d1 + y_0_d2;
  /* fplog32.vhdl:1837:27  */
  assign n4158 = {39'b0, cin_0_d3};  //  uext
  /* fplog32.vhdl:1837:27  */
  assign n4159 = n4157 + n4158;
  /* fplog32.vhdl:1838:14  */
  assign n4160 = s_0[38:0]; // extract
  /* fplog32.vhdl:1839:16  */
  assign n4161 = s_0[39]; // extract
  /* fplog32.vhdl:1840:18  */
  assign n4162 = x[39]; // extract
  /* fplog32.vhdl:1840:15  */
  assign n4164 = {1'b0, n4162};
  /* fplog32.vhdl:1841:18  */
  assign n4165 = y[39]; // extract
  /* fplog32.vhdl:1841:15  */
  assign n4167 = {1'b0, n4165};
  /* fplog32.vhdl:1842:18  */
  assign n4168 = x_1_d1 + y_1_d2;
  /* fplog32.vhdl:1842:27  */
  assign n4169 = {1'b0, cin_1};  //  uext
  /* fplog32.vhdl:1842:27  */
  assign n4170 = n4168 + n4169;
  /* fplog32.vhdl:1843:14  */
  assign n4171 = s_1[0]; // extract
  /* fplog32.vhdl:1844:13  */
  assign n4172 = {r_1, r_0};
  /* fplog32.vhdl:1822:10  */
  always @(posedge clk)
    n4173 <= cin_0;
  /* fplog32.vhdl:1822:10  */
  always @(posedge clk)
    n4174 <= cin_0_d1;
  /* fplog32.vhdl:1822:10  */
  always @(posedge clk)
    n4175 <= cin_0_d2;
  /* fplog32.vhdl:1822:10  */
  always @(posedge clk)
    n4176 <= x_0;
  /* fplog32.vhdl:1822:10  */
  always @(posedge clk)
    n4177 <= y_0;
  /* fplog32.vhdl:1822:10  */
  always @(posedge clk)
    n4178 <= y_0_d1;
  /* fplog32.vhdl:1822:10  */
  always @(posedge clk)
    n4179 <= x_1;
  /* fplog32.vhdl:1822:10  */
  always @(posedge clk)
    n4180 <= y_1;
  /* fplog32.vhdl:1822:10  */
  always @(posedge clk)
    n4181 <= y_1_d1;
endmodule

module logtable1_freq500_uid22
  (input  [6:0] x,
   output [32:0] y);
  wire [32:0] y0;
  wire [32:0] y1;
  wire n3752;
  wire n3755;
  wire n3758;
  wire n3761;
  wire n3764;
  wire n3767;
  wire n3770;
  wire n3773;
  wire n3776;
  wire n3779;
  wire n3782;
  wire n3785;
  wire n3788;
  wire n3791;
  wire n3794;
  wire n3797;
  wire n3800;
  wire n3803;
  wire n3806;
  wire n3809;
  wire n3812;
  wire n3815;
  wire n3818;
  wire n3821;
  wire n3824;
  wire n3827;
  wire n3830;
  wire n3833;
  wire n3836;
  wire n3839;
  wire n3842;
  wire n3845;
  wire n3848;
  wire n3851;
  wire n3854;
  wire n3857;
  wire n3860;
  wire n3863;
  wire n3866;
  wire n3869;
  wire n3872;
  wire n3875;
  wire n3878;
  wire n3881;
  wire n3884;
  wire n3887;
  wire n3890;
  wire n3893;
  wire n3896;
  wire n3899;
  wire n3902;
  wire n3905;
  wire n3908;
  wire n3911;
  wire n3914;
  wire n3917;
  wire n3920;
  wire n3923;
  wire n3926;
  wire n3929;
  wire n3932;
  wire n3935;
  wire n3938;
  wire n3941;
  wire n3944;
  wire n3947;
  wire n3950;
  wire n3953;
  wire n3956;
  wire n3959;
  wire n3962;
  wire n3965;
  wire n3968;
  wire n3971;
  wire n3974;
  wire n3977;
  wire n3980;
  wire n3983;
  wire n3986;
  wire n3989;
  wire n3992;
  wire n3995;
  wire n3998;
  wire n4001;
  wire n4004;
  wire n4007;
  wire n4010;
  wire n4013;
  wire n4016;
  wire n4019;
  wire n4022;
  wire n4025;
  wire n4028;
  wire n4031;
  wire n4034;
  wire n4037;
  wire n4040;
  wire n4043;
  wire n4046;
  wire n4049;
  wire n4052;
  wire n4055;
  wire n4058;
  wire n4061;
  wire n4064;
  wire n4067;
  wire n4070;
  wire n4073;
  wire n4076;
  wire n4079;
  wire n4082;
  wire n4085;
  wire n4088;
  wire n4091;
  wire n4094;
  wire n4097;
  wire n4100;
  wire n4103;
  wire n4106;
  wire n4109;
  wire n4112;
  wire n4115;
  wire n4118;
  wire n4121;
  wire n4124;
  wire n4127;
  wire n4130;
  wire n4133;
  wire [127:0] n4135;
  reg [32:0] n4136;
  assign y = y1; //(module output)
  /* fplog32.vhdl:582:8  */
  assign y0 = n4136; // (signal)
  /* fplog32.vhdl:584:8  */
  assign y1 = y0; // (signal)
  /* fplog32.vhdl:588:43  */
  assign n3752 = x == 7'b0000000;
  /* fplog32.vhdl:589:43  */
  assign n3755 = x == 7'b0000001;
  /* fplog32.vhdl:590:43  */
  assign n3758 = x == 7'b0000010;
  /* fplog32.vhdl:591:43  */
  assign n3761 = x == 7'b0000011;
  /* fplog32.vhdl:592:43  */
  assign n3764 = x == 7'b0000100;
  /* fplog32.vhdl:593:43  */
  assign n3767 = x == 7'b0000101;
  /* fplog32.vhdl:594:43  */
  assign n3770 = x == 7'b0000110;
  /* fplog32.vhdl:595:43  */
  assign n3773 = x == 7'b0000111;
  /* fplog32.vhdl:596:43  */
  assign n3776 = x == 7'b0001000;
  /* fplog32.vhdl:597:43  */
  assign n3779 = x == 7'b0001001;
  /* fplog32.vhdl:598:43  */
  assign n3782 = x == 7'b0001010;
  /* fplog32.vhdl:599:43  */
  assign n3785 = x == 7'b0001011;
  /* fplog32.vhdl:600:43  */
  assign n3788 = x == 7'b0001100;
  /* fplog32.vhdl:601:43  */
  assign n3791 = x == 7'b0001101;
  /* fplog32.vhdl:602:43  */
  assign n3794 = x == 7'b0001110;
  /* fplog32.vhdl:603:43  */
  assign n3797 = x == 7'b0001111;
  /* fplog32.vhdl:604:43  */
  assign n3800 = x == 7'b0010000;
  /* fplog32.vhdl:605:43  */
  assign n3803 = x == 7'b0010001;
  /* fplog32.vhdl:606:43  */
  assign n3806 = x == 7'b0010010;
  /* fplog32.vhdl:607:43  */
  assign n3809 = x == 7'b0010011;
  /* fplog32.vhdl:608:43  */
  assign n3812 = x == 7'b0010100;
  /* fplog32.vhdl:609:43  */
  assign n3815 = x == 7'b0010101;
  /* fplog32.vhdl:610:43  */
  assign n3818 = x == 7'b0010110;
  /* fplog32.vhdl:611:43  */
  assign n3821 = x == 7'b0010111;
  /* fplog32.vhdl:612:43  */
  assign n3824 = x == 7'b0011000;
  /* fplog32.vhdl:613:43  */
  assign n3827 = x == 7'b0011001;
  /* fplog32.vhdl:614:43  */
  assign n3830 = x == 7'b0011010;
  /* fplog32.vhdl:615:43  */
  assign n3833 = x == 7'b0011011;
  /* fplog32.vhdl:616:43  */
  assign n3836 = x == 7'b0011100;
  /* fplog32.vhdl:617:43  */
  assign n3839 = x == 7'b0011101;
  /* fplog32.vhdl:618:43  */
  assign n3842 = x == 7'b0011110;
  /* fplog32.vhdl:619:43  */
  assign n3845 = x == 7'b0011111;
  /* fplog32.vhdl:620:43  */
  assign n3848 = x == 7'b0100000;
  /* fplog32.vhdl:621:43  */
  assign n3851 = x == 7'b0100001;
  /* fplog32.vhdl:622:43  */
  assign n3854 = x == 7'b0100010;
  /* fplog32.vhdl:623:43  */
  assign n3857 = x == 7'b0100011;
  /* fplog32.vhdl:624:43  */
  assign n3860 = x == 7'b0100100;
  /* fplog32.vhdl:625:43  */
  assign n3863 = x == 7'b0100101;
  /* fplog32.vhdl:626:43  */
  assign n3866 = x == 7'b0100110;
  /* fplog32.vhdl:627:43  */
  assign n3869 = x == 7'b0100111;
  /* fplog32.vhdl:628:43  */
  assign n3872 = x == 7'b0101000;
  /* fplog32.vhdl:629:43  */
  assign n3875 = x == 7'b0101001;
  /* fplog32.vhdl:630:43  */
  assign n3878 = x == 7'b0101010;
  /* fplog32.vhdl:631:43  */
  assign n3881 = x == 7'b0101011;
  /* fplog32.vhdl:632:43  */
  assign n3884 = x == 7'b0101100;
  /* fplog32.vhdl:633:43  */
  assign n3887 = x == 7'b0101101;
  /* fplog32.vhdl:634:43  */
  assign n3890 = x == 7'b0101110;
  /* fplog32.vhdl:635:43  */
  assign n3893 = x == 7'b0101111;
  /* fplog32.vhdl:636:43  */
  assign n3896 = x == 7'b0110000;
  /* fplog32.vhdl:637:43  */
  assign n3899 = x == 7'b0110001;
  /* fplog32.vhdl:638:43  */
  assign n3902 = x == 7'b0110010;
  /* fplog32.vhdl:639:43  */
  assign n3905 = x == 7'b0110011;
  /* fplog32.vhdl:640:43  */
  assign n3908 = x == 7'b0110100;
  /* fplog32.vhdl:641:43  */
  assign n3911 = x == 7'b0110101;
  /* fplog32.vhdl:642:43  */
  assign n3914 = x == 7'b0110110;
  /* fplog32.vhdl:643:43  */
  assign n3917 = x == 7'b0110111;
  /* fplog32.vhdl:644:43  */
  assign n3920 = x == 7'b0111000;
  /* fplog32.vhdl:645:43  */
  assign n3923 = x == 7'b0111001;
  /* fplog32.vhdl:646:43  */
  assign n3926 = x == 7'b0111010;
  /* fplog32.vhdl:647:43  */
  assign n3929 = x == 7'b0111011;
  /* fplog32.vhdl:648:43  */
  assign n3932 = x == 7'b0111100;
  /* fplog32.vhdl:649:43  */
  assign n3935 = x == 7'b0111101;
  /* fplog32.vhdl:650:43  */
  assign n3938 = x == 7'b0111110;
  /* fplog32.vhdl:651:43  */
  assign n3941 = x == 7'b0111111;
  /* fplog32.vhdl:652:43  */
  assign n3944 = x == 7'b1000000;
  /* fplog32.vhdl:653:43  */
  assign n3947 = x == 7'b1000001;
  /* fplog32.vhdl:654:43  */
  assign n3950 = x == 7'b1000010;
  /* fplog32.vhdl:655:43  */
  assign n3953 = x == 7'b1000011;
  /* fplog32.vhdl:656:43  */
  assign n3956 = x == 7'b1000100;
  /* fplog32.vhdl:657:43  */
  assign n3959 = x == 7'b1000101;
  /* fplog32.vhdl:658:43  */
  assign n3962 = x == 7'b1000110;
  /* fplog32.vhdl:659:43  */
  assign n3965 = x == 7'b1000111;
  /* fplog32.vhdl:660:43  */
  assign n3968 = x == 7'b1001000;
  /* fplog32.vhdl:661:43  */
  assign n3971 = x == 7'b1001001;
  /* fplog32.vhdl:662:43  */
  assign n3974 = x == 7'b1001010;
  /* fplog32.vhdl:663:43  */
  assign n3977 = x == 7'b1001011;
  /* fplog32.vhdl:664:43  */
  assign n3980 = x == 7'b1001100;
  /* fplog32.vhdl:665:43  */
  assign n3983 = x == 7'b1001101;
  /* fplog32.vhdl:666:43  */
  assign n3986 = x == 7'b1001110;
  /* fplog32.vhdl:667:43  */
  assign n3989 = x == 7'b1001111;
  /* fplog32.vhdl:668:43  */
  assign n3992 = x == 7'b1010000;
  /* fplog32.vhdl:669:43  */
  assign n3995 = x == 7'b1010001;
  /* fplog32.vhdl:670:43  */
  assign n3998 = x == 7'b1010010;
  /* fplog32.vhdl:671:43  */
  assign n4001 = x == 7'b1010011;
  /* fplog32.vhdl:672:43  */
  assign n4004 = x == 7'b1010100;
  /* fplog32.vhdl:673:43  */
  assign n4007 = x == 7'b1010101;
  /* fplog32.vhdl:674:43  */
  assign n4010 = x == 7'b1010110;
  /* fplog32.vhdl:675:43  */
  assign n4013 = x == 7'b1010111;
  /* fplog32.vhdl:676:43  */
  assign n4016 = x == 7'b1011000;
  /* fplog32.vhdl:677:43  */
  assign n4019 = x == 7'b1011001;
  /* fplog32.vhdl:678:43  */
  assign n4022 = x == 7'b1011010;
  /* fplog32.vhdl:679:43  */
  assign n4025 = x == 7'b1011011;
  /* fplog32.vhdl:680:43  */
  assign n4028 = x == 7'b1011100;
  /* fplog32.vhdl:681:43  */
  assign n4031 = x == 7'b1011101;
  /* fplog32.vhdl:682:43  */
  assign n4034 = x == 7'b1011110;
  /* fplog32.vhdl:683:43  */
  assign n4037 = x == 7'b1011111;
  /* fplog32.vhdl:684:43  */
  assign n4040 = x == 7'b1100000;
  /* fplog32.vhdl:685:43  */
  assign n4043 = x == 7'b1100001;
  /* fplog32.vhdl:686:43  */
  assign n4046 = x == 7'b1100010;
  /* fplog32.vhdl:687:43  */
  assign n4049 = x == 7'b1100011;
  /* fplog32.vhdl:688:43  */
  assign n4052 = x == 7'b1100100;
  /* fplog32.vhdl:689:43  */
  assign n4055 = x == 7'b1100101;
  /* fplog32.vhdl:690:43  */
  assign n4058 = x == 7'b1100110;
  /* fplog32.vhdl:691:43  */
  assign n4061 = x == 7'b1100111;
  /* fplog32.vhdl:692:43  */
  assign n4064 = x == 7'b1101000;
  /* fplog32.vhdl:693:43  */
  assign n4067 = x == 7'b1101001;
  /* fplog32.vhdl:694:43  */
  assign n4070 = x == 7'b1101010;
  /* fplog32.vhdl:695:43  */
  assign n4073 = x == 7'b1101011;
  /* fplog32.vhdl:696:43  */
  assign n4076 = x == 7'b1101100;
  /* fplog32.vhdl:697:43  */
  assign n4079 = x == 7'b1101101;
  /* fplog32.vhdl:698:43  */
  assign n4082 = x == 7'b1101110;
  /* fplog32.vhdl:699:43  */
  assign n4085 = x == 7'b1101111;
  /* fplog32.vhdl:700:43  */
  assign n4088 = x == 7'b1110000;
  /* fplog32.vhdl:701:43  */
  assign n4091 = x == 7'b1110001;
  /* fplog32.vhdl:702:43  */
  assign n4094 = x == 7'b1110010;
  /* fplog32.vhdl:703:43  */
  assign n4097 = x == 7'b1110011;
  /* fplog32.vhdl:704:43  */
  assign n4100 = x == 7'b1110100;
  /* fplog32.vhdl:705:43  */
  assign n4103 = x == 7'b1110101;
  /* fplog32.vhdl:706:43  */
  assign n4106 = x == 7'b1110110;
  /* fplog32.vhdl:707:43  */
  assign n4109 = x == 7'b1110111;
  /* fplog32.vhdl:708:43  */
  assign n4112 = x == 7'b1111000;
  /* fplog32.vhdl:709:43  */
  assign n4115 = x == 7'b1111001;
  /* fplog32.vhdl:710:43  */
  assign n4118 = x == 7'b1111010;
  /* fplog32.vhdl:711:43  */
  assign n4121 = x == 7'b1111011;
  /* fplog32.vhdl:712:43  */
  assign n4124 = x == 7'b1111100;
  /* fplog32.vhdl:713:43  */
  assign n4127 = x == 7'b1111101;
  /* fplog32.vhdl:714:43  */
  assign n4130 = x == 7'b1111110;
  /* fplog32.vhdl:715:43  */
  assign n4133 = x == 7'b1111111;
  assign n4135 = {n4133, n4130, n4127, n4124, n4121, n4118, n4115, n4112, n4109, n4106, n4103, n4100, n4097, n4094, n4091, n4088, n4085, n4082, n4079, n4076, n4073, n4070, n4067, n4064, n4061, n4058, n4055, n4052, n4049, n4046, n4043, n4040, n4037, n4034, n4031, n4028, n4025, n4022, n4019, n4016, n4013, n4010, n4007, n4004, n4001, n3998, n3995, n3992, n3989, n3986, n3983, n3980, n3977, n3974, n3971, n3968, n3965, n3962, n3959, n3956, n3953, n3950, n3947, n3944, n3941, n3938, n3935, n3932, n3929, n3926, n3923, n3920, n3917, n3914, n3911, n3908, n3905, n3902, n3899, n3896, n3893, n3890, n3887, n3884, n3881, n3878, n3875, n3872, n3869, n3866, n3863, n3860, n3857, n3854, n3851, n3848, n3845, n3842, n3839, n3836, n3833, n3830, n3827, n3824, n3821, n3818, n3815, n3812, n3809, n3806, n3803, n3800, n3797, n3794, n3791, n3788, n3785, n3782, n3779, n3776, n3773, n3770, n3767, n3764, n3761, n3758, n3755, n3752};
  /* fplog32.vhdl:587:4  */
  always @*
    case (n4135)
      128'b10000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n4136 = 33'b111111101111100101010111011110001;
      128'b01000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n4136 = 33'b111111001111010101100011101110001;
      128'b00100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n4136 = 33'b111110101111000101111000000110001;
      128'b00010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n4136 = 33'b111110001110110110010100100101111;
      128'b00001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n4136 = 33'b111101101110100110111001001101011;
      128'b00000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n4136 = 33'b111101001110010111100101111100101;
      128'b00000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n4136 = 33'b111100101110001000011010110011100;
      128'b00000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n4136 = 33'b111100001101111001010111110001111;
      128'b00000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n4136 = 33'b111011101101101010011100110111111;
      128'b00000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n4136 = 33'b111011001101011011101010000101011;
      128'b00000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n4136 = 33'b111010101101001100111111011010001;
      128'b00000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n4136 = 33'b111010001100111110011100110110011;
      128'b00000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n4136 = 33'b111001101100110000000010011001110;
      128'b00000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n4136 = 33'b111001001100100001110000000100011;
      128'b00000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n4136 = 33'b111000101100010011100101110110001;
      128'b00000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n4136 = 33'b111000001100000101100011101111000;
      128'b00000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n4136 = 33'b110111101011110111101001101110110;
      128'b00000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n4136 = 33'b110111001011101001110111110101100;
      128'b00000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n4136 = 33'b110110101011011100001110000011010;
      128'b00000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n4136 = 33'b110110001011001110101100010111110;
      128'b00000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n4136 = 33'b110101101011000001010010110010111;
      128'b00000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n4136 = 33'b110101001010110100000001010100111;
      128'b00000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n4136 = 33'b110100101010100110110111111101011;
      128'b00000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n4136 = 33'b110100001010011001110110101100100;
      128'b00000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n4136 = 33'b110011101010001100111101100010001;
      128'b00000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n4136 = 33'b110011001010000000001100011110001;
      128'b00000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n4136 = 33'b110010101001110011100011100000101;
      128'b00000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n4136 = 33'b110010001001100111000010101001010;
      128'b00000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n4136 = 33'b110001101001011010101001111000010;
      128'b00000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n4136 = 33'b110001001001001110011001001101011;
      128'b00000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n4136 = 33'b110000101001000010010000101000110;
      128'b00000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n4136 = 33'b110000001000110110010000001010000;
      128'b00000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n4136 = 33'b101111101000101010010111110001011;
      128'b00000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n4136 = 33'b101111001000011110100111011110100;
      128'b00000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n4136 = 33'b101110101000010010111111010001101;
      128'b00000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n4136 = 33'b101110001000000111011111001010100;
      128'b00000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n4136 = 33'b101101100111111100000111001001001;
      128'b00000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n4136 = 33'b101101000111110000110111001101100;
      128'b00000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n4136 = 33'b101100100111100101101111010111011;
      128'b00000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n4136 = 33'b101100000111011010101111100110111;
      128'b00000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n4136 = 33'b101011100111001111110111111011110;
      128'b00000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n4136 = 33'b101011000111000101001000010110001;
      128'b00000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n4136 = 33'b101010100110111010100000110101111;
      128'b00000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n4136 = 33'b101010000110110000000001011010111;
      128'b00000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000: n4136 = 33'b101001100110100101101010000101000;
      128'b00000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000: n4136 = 33'b101001000110011011011010110100100;
      128'b00000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000: n4136 = 33'b101000100110010001010011101001000;
      128'b00000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000: n4136 = 33'b101000000110000111010100100010100;
      128'b00000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000: n4136 = 33'b100111100101111101011101100001000;
      128'b00000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000: n4136 = 33'b100111000101110011101110100100011;
      128'b00000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000: n4136 = 33'b100110100101101010000111101100101;
      128'b00000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000: n4136 = 33'b100110000101100000101000111001101;
      128'b00000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000: n4136 = 33'b100101100101010111010010001011011;
      128'b00000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000: n4136 = 33'b100101000101001110000011100001111;
      128'b00000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000: n4136 = 33'b100100100101000100111100111100111;
      128'b00000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000: n4136 = 33'b100100000100111011111110011100011;
      128'b00000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000: n4136 = 33'b100011100100110011001000000000011;
      128'b00000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000: n4136 = 33'b100011000100101010011001101000111;
      128'b00000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000: n4136 = 33'b100010100100100001110011010101101;
      128'b00000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000: n4136 = 33'b100010000100011001010101000110101;
      128'b00000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000: n4136 = 33'b100001100100010000111110111011111;
      128'b00000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000: n4136 = 33'b100001000100001000110000110101010;
      128'b00000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000: n4136 = 33'b100000100100000000101010110010110;
      128'b00000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000: n4136 = 33'b100000000011111000101100110100010;
      128'b00000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000: n4136 = 33'b011111110011110100110000110110100;
      128'b00000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000: n4136 = 33'b011111010011101100111110111101111;
      128'b00000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000: n4136 = 33'b011110110011100101010101001001001;
      128'b00000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000: n4136 = 33'b011110010011011101110011011000010;
      128'b00000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000: n4136 = 33'b011101110011010110011001101011000;
      128'b00000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000: n4136 = 33'b011101010011001111001000000001100;
      128'b00000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000: n4136 = 33'b011100110011000111111110011011101;
      128'b00000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000: n4136 = 33'b011100010011000000111100111001010;
      128'b00000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000: n4136 = 33'b011011110010111010000011011010100;
      128'b00000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000: n4136 = 33'b011011010010110011010001111111000;
      128'b00000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000: n4136 = 33'b011010110010101100101000100111000;
      128'b00000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000: n4136 = 33'b011010010010100110000111010010010;
      128'b00000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000: n4136 = 33'b011001110010011111101110000000101;
      128'b00000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000: n4136 = 33'b011001010010011001011100110010010;
      128'b00000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000: n4136 = 33'b011000110010010011010011100111000;
      128'b00000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000: n4136 = 33'b011000010010001101010010011110110;
      128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000: n4136 = 33'b010111110010000111011001011001100;
      128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000: n4136 = 33'b010111010010000001101000010111010;
      128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000: n4136 = 33'b010110110001111011111111010111110;
      128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000: n4136 = 33'b010110010001110110011110011011001;
      128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000: n4136 = 33'b010101110001110001000101100001010;
      128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000: n4136 = 33'b010101010001101011110100101010000;
      128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000: n4136 = 33'b010100110001100110101011110101010;
      128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000: n4136 = 33'b010100010001100001101011000011001;
      128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000: n4136 = 33'b010011110001011100110010010011100;
      128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000: n4136 = 33'b010011010001011000000001100110010;
      128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000: n4136 = 33'b010010110001010011011000111011011;
      128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000: n4136 = 33'b010010010001001110111000010010110;
      128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000: n4136 = 33'b010001110001001010011111101100100;
      128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000: n4136 = 33'b010001010001000110001111001000010;
      128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000: n4136 = 33'b010000110001000010000110100110001;
      128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000: n4136 = 33'b010000010000111110000110000110000;
      128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000: n4136 = 33'b001111110000111010001101101000000;
      128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000: n4136 = 33'b001111010000110110011101001011110;
      128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000: n4136 = 33'b001110110000110010110100110001100;
      128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000: n4136 = 33'b001110010000101111010100011000111;
      128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000: n4136 = 33'b001101110000101011111100000010001;
      128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000: n4136 = 33'b001101010000101000101011101101000;
      128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000: n4136 = 33'b001100110000100101100011011001011;
      128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000: n4136 = 33'b001100010000100010100011000111011;
      128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000: n4136 = 33'b001011110000011111101010110110110;
      128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000: n4136 = 33'b001011010000011100111010100111101;
      128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000: n4136 = 33'b001010110000011010010010011001110;
      128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000: n4136 = 33'b001010010000010111110010001101010;
      128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000: n4136 = 33'b001001110000010101011010000010000;
      128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000: n4136 = 33'b001001010000010011001001110111111;
      128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000: n4136 = 33'b001000110000010001000001101110111;
      128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000: n4136 = 33'b001000010000001111000001100110110;
      128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000: n4136 = 33'b000111110000001101001001011111110;
      128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000: n4136 = 33'b000111010000001011011001011001101;
      128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000: n4136 = 33'b000110110000001001110001010100011;
      128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000: n4136 = 33'b000110010000001000010001001111111;
      128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000: n4136 = 33'b000101110000000110111001001100000;
      128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000: n4136 = 33'b000101010000000101101001001001000;
      128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000: n4136 = 33'b000100110000000100100001000110011;
      128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000: n4136 = 33'b000100010000000011100001000100011;
      128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000: n4136 = 33'b000011110000000010101001000010111;
      128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000: n4136 = 33'b000011010000000001111001000001110;
      128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000: n4136 = 33'b000010110000000001010001000001000;
      128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000: n4136 = 33'b000010010000000000110001000000100;
      128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000: n4136 = 33'b000001110000000000011001000000001;
      128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100: n4136 = 33'b000001010000000000001001000000000;
      128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010: n4136 = 33'b000000110000000000000001000000000;
      128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001: n4136 = 33'b000000010000000000000001000000000;
      default: n4136 = 33'bX;
    endcase
endmodule

module logtable0_freq500_uid20
  (input  clk,
   input  [8:0] x,
   output [39:0] y);
  wire [39:0] y0;
  wire [39:0] y0_d1;
  wire [39:0] y1;
  wire [8:0] x_d1;
  wire n2210;
  wire n2213;
  wire n2216;
  wire n2219;
  wire n2222;
  wire n2225;
  wire n2228;
  wire n2231;
  wire n2234;
  wire n2237;
  wire n2240;
  wire n2243;
  wire n2246;
  wire n2249;
  wire n2252;
  wire n2255;
  wire n2258;
  wire n2261;
  wire n2264;
  wire n2267;
  wire n2270;
  wire n2273;
  wire n2276;
  wire n2279;
  wire n2282;
  wire n2285;
  wire n2288;
  wire n2291;
  wire n2294;
  wire n2297;
  wire n2300;
  wire n2303;
  wire n2306;
  wire n2309;
  wire n2312;
  wire n2315;
  wire n2318;
  wire n2321;
  wire n2324;
  wire n2327;
  wire n2330;
  wire n2333;
  wire n2336;
  wire n2339;
  wire n2342;
  wire n2345;
  wire n2348;
  wire n2351;
  wire n2354;
  wire n2357;
  wire n2360;
  wire n2363;
  wire n2366;
  wire n2369;
  wire n2372;
  wire n2375;
  wire n2378;
  wire n2381;
  wire n2384;
  wire n2387;
  wire n2390;
  wire n2393;
  wire n2396;
  wire n2399;
  wire n2402;
  wire n2405;
  wire n2408;
  wire n2411;
  wire n2414;
  wire n2417;
  wire n2420;
  wire n2423;
  wire n2426;
  wire n2429;
  wire n2432;
  wire n2435;
  wire n2438;
  wire n2441;
  wire n2444;
  wire n2447;
  wire n2450;
  wire n2453;
  wire n2456;
  wire n2459;
  wire n2462;
  wire n2465;
  wire n2468;
  wire n2471;
  wire n2474;
  wire n2477;
  wire n2480;
  wire n2483;
  wire n2486;
  wire n2489;
  wire n2492;
  wire n2495;
  wire n2498;
  wire n2501;
  wire n2504;
  wire n2507;
  wire n2510;
  wire n2513;
  wire n2516;
  wire n2519;
  wire n2522;
  wire n2525;
  wire n2528;
  wire n2531;
  wire n2534;
  wire n2537;
  wire n2540;
  wire n2543;
  wire n2546;
  wire n2549;
  wire n2552;
  wire n2555;
  wire n2558;
  wire n2561;
  wire n2564;
  wire n2567;
  wire n2570;
  wire n2573;
  wire n2576;
  wire n2579;
  wire n2582;
  wire n2585;
  wire n2588;
  wire n2591;
  wire n2594;
  wire n2597;
  wire n2600;
  wire n2603;
  wire n2606;
  wire n2609;
  wire n2612;
  wire n2615;
  wire n2618;
  wire n2621;
  wire n2624;
  wire n2627;
  wire n2630;
  wire n2633;
  wire n2636;
  wire n2639;
  wire n2642;
  wire n2645;
  wire n2648;
  wire n2651;
  wire n2654;
  wire n2657;
  wire n2660;
  wire n2663;
  wire n2666;
  wire n2669;
  wire n2672;
  wire n2675;
  wire n2678;
  wire n2681;
  wire n2684;
  wire n2687;
  wire n2690;
  wire n2693;
  wire n2696;
  wire n2699;
  wire n2702;
  wire n2705;
  wire n2708;
  wire n2711;
  wire n2714;
  wire n2717;
  wire n2720;
  wire n2723;
  wire n2726;
  wire n2729;
  wire n2732;
  wire n2735;
  wire n2738;
  wire n2741;
  wire n2744;
  wire n2747;
  wire n2750;
  wire n2753;
  wire n2756;
  wire n2759;
  wire n2762;
  wire n2765;
  wire n2768;
  wire n2771;
  wire n2774;
  wire n2777;
  wire n2780;
  wire n2783;
  wire n2786;
  wire n2789;
  wire n2792;
  wire n2795;
  wire n2798;
  wire n2801;
  wire n2804;
  wire n2807;
  wire n2810;
  wire n2813;
  wire n2816;
  wire n2819;
  wire n2822;
  wire n2825;
  wire n2828;
  wire n2831;
  wire n2834;
  wire n2837;
  wire n2840;
  wire n2843;
  wire n2846;
  wire n2849;
  wire n2852;
  wire n2855;
  wire n2858;
  wire n2861;
  wire n2864;
  wire n2867;
  wire n2870;
  wire n2873;
  wire n2876;
  wire n2879;
  wire n2882;
  wire n2885;
  wire n2888;
  wire n2891;
  wire n2894;
  wire n2897;
  wire n2900;
  wire n2903;
  wire n2906;
  wire n2909;
  wire n2912;
  wire n2915;
  wire n2918;
  wire n2921;
  wire n2924;
  wire n2927;
  wire n2930;
  wire n2933;
  wire n2936;
  wire n2939;
  wire n2942;
  wire n2945;
  wire n2948;
  wire n2951;
  wire n2954;
  wire n2957;
  wire n2960;
  wire n2963;
  wire n2966;
  wire n2969;
  wire n2972;
  wire n2975;
  wire n2978;
  wire n2981;
  wire n2984;
  wire n2987;
  wire n2990;
  wire n2993;
  wire n2996;
  wire n2999;
  wire n3002;
  wire n3005;
  wire n3008;
  wire n3011;
  wire n3014;
  wire n3017;
  wire n3020;
  wire n3023;
  wire n3026;
  wire n3029;
  wire n3032;
  wire n3035;
  wire n3038;
  wire n3041;
  wire n3044;
  wire n3047;
  wire n3050;
  wire n3053;
  wire n3056;
  wire n3059;
  wire n3062;
  wire n3065;
  wire n3068;
  wire n3071;
  wire n3074;
  wire n3077;
  wire n3080;
  wire n3083;
  wire n3086;
  wire n3089;
  wire n3092;
  wire n3095;
  wire n3098;
  wire n3101;
  wire n3104;
  wire n3107;
  wire n3110;
  wire n3113;
  wire n3116;
  wire n3119;
  wire n3122;
  wire n3125;
  wire n3128;
  wire n3131;
  wire n3134;
  wire n3137;
  wire n3140;
  wire n3143;
  wire n3146;
  wire n3149;
  wire n3152;
  wire n3155;
  wire n3158;
  wire n3161;
  wire n3164;
  wire n3167;
  wire n3170;
  wire n3173;
  wire n3176;
  wire n3179;
  wire n3182;
  wire n3185;
  wire n3188;
  wire n3191;
  wire n3194;
  wire n3197;
  wire n3200;
  wire n3203;
  wire n3206;
  wire n3209;
  wire n3212;
  wire n3215;
  wire n3218;
  wire n3221;
  wire n3224;
  wire n3227;
  wire n3230;
  wire n3233;
  wire n3236;
  wire n3239;
  wire n3242;
  wire n3245;
  wire n3248;
  wire n3251;
  wire n3254;
  wire n3257;
  wire n3260;
  wire n3263;
  wire n3266;
  wire n3269;
  wire n3272;
  wire n3275;
  wire n3278;
  wire n3281;
  wire n3284;
  wire n3287;
  wire n3290;
  wire n3293;
  wire n3296;
  wire n3299;
  wire n3302;
  wire n3305;
  wire n3308;
  wire n3311;
  wire n3314;
  wire n3317;
  wire n3320;
  wire n3323;
  wire n3326;
  wire n3329;
  wire n3332;
  wire n3335;
  wire n3338;
  wire n3341;
  wire n3344;
  wire n3347;
  wire n3350;
  wire n3353;
  wire n3356;
  wire n3359;
  wire n3362;
  wire n3365;
  wire n3368;
  wire n3371;
  wire n3374;
  wire n3377;
  wire n3380;
  wire n3383;
  wire n3386;
  wire n3389;
  wire n3392;
  wire n3395;
  wire n3398;
  wire n3401;
  wire n3404;
  wire n3407;
  wire n3410;
  wire n3413;
  wire n3416;
  wire n3419;
  wire n3422;
  wire n3425;
  wire n3428;
  wire n3431;
  wire n3434;
  wire n3437;
  wire n3440;
  wire n3443;
  wire n3446;
  wire n3449;
  wire n3452;
  wire n3455;
  wire n3458;
  wire n3461;
  wire n3464;
  wire n3467;
  wire n3470;
  wire n3473;
  wire n3476;
  wire n3479;
  wire n3482;
  wire n3485;
  wire n3488;
  wire n3491;
  wire n3494;
  wire n3497;
  wire n3500;
  wire n3503;
  wire n3506;
  wire n3509;
  wire n3512;
  wire n3515;
  wire n3518;
  wire n3521;
  wire n3524;
  wire n3527;
  wire n3530;
  wire n3533;
  wire n3536;
  wire n3539;
  wire n3542;
  wire n3545;
  wire n3548;
  wire n3551;
  wire n3554;
  wire n3557;
  wire n3560;
  wire n3563;
  wire n3566;
  wire n3569;
  wire n3572;
  wire n3575;
  wire n3578;
  wire n3581;
  wire n3584;
  wire n3587;
  wire n3590;
  wire n3593;
  wire n3596;
  wire n3599;
  wire n3602;
  wire n3605;
  wire n3608;
  wire n3611;
  wire n3614;
  wire n3617;
  wire n3620;
  wire n3623;
  wire n3626;
  wire n3629;
  wire n3632;
  wire n3635;
  wire n3638;
  wire n3641;
  wire n3644;
  wire n3647;
  wire n3650;
  wire n3653;
  wire n3656;
  wire n3659;
  wire n3662;
  wire n3665;
  wire n3668;
  wire n3671;
  wire n3674;
  wire n3677;
  wire n3680;
  wire n3683;
  wire n3686;
  wire n3689;
  wire n3692;
  wire n3695;
  wire n3698;
  wire n3701;
  wire n3704;
  wire n3707;
  wire n3710;
  wire n3713;
  wire n3716;
  wire n3719;
  wire n3722;
  wire n3725;
  wire n3728;
  wire n3731;
  wire n3734;
  wire n3737;
  wire n3740;
  wire n3743;
  wire [511:0] n3745;
  reg [39:0] n3746;
  reg [39:0] n3747;
  reg [8:0] n3748;
  assign y = y1; //(module output)
  /* fplog32.vhdl:1235:8  */
  assign y0 = n3746; // (signal)
  /* fplog32.vhdl:1235:12  */
  assign y0_d1 = n3747; // (signal)
  /* fplog32.vhdl:1237:8  */
  assign y1 = y0_d1; // (signal)
  /* fplog32.vhdl:1239:8  */
  assign x_d1 = n3748; // (signal)
  /* fplog32.vhdl:1250:50  */
  assign n2210 = x_d1 == 9'b000000000;
  /* fplog32.vhdl:1251:50  */
  assign n2213 = x_d1 == 9'b000000001;
  /* fplog32.vhdl:1252:50  */
  assign n2216 = x_d1 == 9'b000000010;
  /* fplog32.vhdl:1253:50  */
  assign n2219 = x_d1 == 9'b000000011;
  /* fplog32.vhdl:1254:50  */
  assign n2222 = x_d1 == 9'b000000100;
  /* fplog32.vhdl:1255:50  */
  assign n2225 = x_d1 == 9'b000000101;
  /* fplog32.vhdl:1256:50  */
  assign n2228 = x_d1 == 9'b000000110;
  /* fplog32.vhdl:1257:50  */
  assign n2231 = x_d1 == 9'b000000111;
  /* fplog32.vhdl:1258:50  */
  assign n2234 = x_d1 == 9'b000001000;
  /* fplog32.vhdl:1259:50  */
  assign n2237 = x_d1 == 9'b000001001;
  /* fplog32.vhdl:1260:50  */
  assign n2240 = x_d1 == 9'b000001010;
  /* fplog32.vhdl:1261:50  */
  assign n2243 = x_d1 == 9'b000001011;
  /* fplog32.vhdl:1262:50  */
  assign n2246 = x_d1 == 9'b000001100;
  /* fplog32.vhdl:1263:50  */
  assign n2249 = x_d1 == 9'b000001101;
  /* fplog32.vhdl:1264:50  */
  assign n2252 = x_d1 == 9'b000001110;
  /* fplog32.vhdl:1265:50  */
  assign n2255 = x_d1 == 9'b000001111;
  /* fplog32.vhdl:1266:50  */
  assign n2258 = x_d1 == 9'b000010000;
  /* fplog32.vhdl:1267:50  */
  assign n2261 = x_d1 == 9'b000010001;
  /* fplog32.vhdl:1268:50  */
  assign n2264 = x_d1 == 9'b000010010;
  /* fplog32.vhdl:1269:50  */
  assign n2267 = x_d1 == 9'b000010011;
  /* fplog32.vhdl:1270:50  */
  assign n2270 = x_d1 == 9'b000010100;
  /* fplog32.vhdl:1271:50  */
  assign n2273 = x_d1 == 9'b000010101;
  /* fplog32.vhdl:1272:50  */
  assign n2276 = x_d1 == 9'b000010110;
  /* fplog32.vhdl:1273:50  */
  assign n2279 = x_d1 == 9'b000010111;
  /* fplog32.vhdl:1274:50  */
  assign n2282 = x_d1 == 9'b000011000;
  /* fplog32.vhdl:1275:50  */
  assign n2285 = x_d1 == 9'b000011001;
  /* fplog32.vhdl:1276:50  */
  assign n2288 = x_d1 == 9'b000011010;
  /* fplog32.vhdl:1277:50  */
  assign n2291 = x_d1 == 9'b000011011;
  /* fplog32.vhdl:1278:50  */
  assign n2294 = x_d1 == 9'b000011100;
  /* fplog32.vhdl:1279:50  */
  assign n2297 = x_d1 == 9'b000011101;
  /* fplog32.vhdl:1280:50  */
  assign n2300 = x_d1 == 9'b000011110;
  /* fplog32.vhdl:1281:50  */
  assign n2303 = x_d1 == 9'b000011111;
  /* fplog32.vhdl:1282:50  */
  assign n2306 = x_d1 == 9'b000100000;
  /* fplog32.vhdl:1283:50  */
  assign n2309 = x_d1 == 9'b000100001;
  /* fplog32.vhdl:1284:50  */
  assign n2312 = x_d1 == 9'b000100010;
  /* fplog32.vhdl:1285:50  */
  assign n2315 = x_d1 == 9'b000100011;
  /* fplog32.vhdl:1286:50  */
  assign n2318 = x_d1 == 9'b000100100;
  /* fplog32.vhdl:1287:50  */
  assign n2321 = x_d1 == 9'b000100101;
  /* fplog32.vhdl:1288:50  */
  assign n2324 = x_d1 == 9'b000100110;
  /* fplog32.vhdl:1289:50  */
  assign n2327 = x_d1 == 9'b000100111;
  /* fplog32.vhdl:1290:50  */
  assign n2330 = x_d1 == 9'b000101000;
  /* fplog32.vhdl:1291:50  */
  assign n2333 = x_d1 == 9'b000101001;
  /* fplog32.vhdl:1292:50  */
  assign n2336 = x_d1 == 9'b000101010;
  /* fplog32.vhdl:1293:50  */
  assign n2339 = x_d1 == 9'b000101011;
  /* fplog32.vhdl:1294:50  */
  assign n2342 = x_d1 == 9'b000101100;
  /* fplog32.vhdl:1295:50  */
  assign n2345 = x_d1 == 9'b000101101;
  /* fplog32.vhdl:1296:50  */
  assign n2348 = x_d1 == 9'b000101110;
  /* fplog32.vhdl:1297:50  */
  assign n2351 = x_d1 == 9'b000101111;
  /* fplog32.vhdl:1298:50  */
  assign n2354 = x_d1 == 9'b000110000;
  /* fplog32.vhdl:1299:50  */
  assign n2357 = x_d1 == 9'b000110001;
  /* fplog32.vhdl:1300:50  */
  assign n2360 = x_d1 == 9'b000110010;
  /* fplog32.vhdl:1301:50  */
  assign n2363 = x_d1 == 9'b000110011;
  /* fplog32.vhdl:1302:50  */
  assign n2366 = x_d1 == 9'b000110100;
  /* fplog32.vhdl:1303:50  */
  assign n2369 = x_d1 == 9'b000110101;
  /* fplog32.vhdl:1304:50  */
  assign n2372 = x_d1 == 9'b000110110;
  /* fplog32.vhdl:1305:50  */
  assign n2375 = x_d1 == 9'b000110111;
  /* fplog32.vhdl:1306:50  */
  assign n2378 = x_d1 == 9'b000111000;
  /* fplog32.vhdl:1307:50  */
  assign n2381 = x_d1 == 9'b000111001;
  /* fplog32.vhdl:1308:50  */
  assign n2384 = x_d1 == 9'b000111010;
  /* fplog32.vhdl:1309:50  */
  assign n2387 = x_d1 == 9'b000111011;
  /* fplog32.vhdl:1310:50  */
  assign n2390 = x_d1 == 9'b000111100;
  /* fplog32.vhdl:1311:50  */
  assign n2393 = x_d1 == 9'b000111101;
  /* fplog32.vhdl:1312:50  */
  assign n2396 = x_d1 == 9'b000111110;
  /* fplog32.vhdl:1313:50  */
  assign n2399 = x_d1 == 9'b000111111;
  /* fplog32.vhdl:1314:50  */
  assign n2402 = x_d1 == 9'b001000000;
  /* fplog32.vhdl:1315:50  */
  assign n2405 = x_d1 == 9'b001000001;
  /* fplog32.vhdl:1316:50  */
  assign n2408 = x_d1 == 9'b001000010;
  /* fplog32.vhdl:1317:50  */
  assign n2411 = x_d1 == 9'b001000011;
  /* fplog32.vhdl:1318:50  */
  assign n2414 = x_d1 == 9'b001000100;
  /* fplog32.vhdl:1319:50  */
  assign n2417 = x_d1 == 9'b001000101;
  /* fplog32.vhdl:1320:50  */
  assign n2420 = x_d1 == 9'b001000110;
  /* fplog32.vhdl:1321:50  */
  assign n2423 = x_d1 == 9'b001000111;
  /* fplog32.vhdl:1322:50  */
  assign n2426 = x_d1 == 9'b001001000;
  /* fplog32.vhdl:1323:50  */
  assign n2429 = x_d1 == 9'b001001001;
  /* fplog32.vhdl:1324:50  */
  assign n2432 = x_d1 == 9'b001001010;
  /* fplog32.vhdl:1325:50  */
  assign n2435 = x_d1 == 9'b001001011;
  /* fplog32.vhdl:1326:50  */
  assign n2438 = x_d1 == 9'b001001100;
  /* fplog32.vhdl:1327:50  */
  assign n2441 = x_d1 == 9'b001001101;
  /* fplog32.vhdl:1328:50  */
  assign n2444 = x_d1 == 9'b001001110;
  /* fplog32.vhdl:1329:50  */
  assign n2447 = x_d1 == 9'b001001111;
  /* fplog32.vhdl:1330:50  */
  assign n2450 = x_d1 == 9'b001010000;
  /* fplog32.vhdl:1331:50  */
  assign n2453 = x_d1 == 9'b001010001;
  /* fplog32.vhdl:1332:50  */
  assign n2456 = x_d1 == 9'b001010010;
  /* fplog32.vhdl:1333:50  */
  assign n2459 = x_d1 == 9'b001010011;
  /* fplog32.vhdl:1334:50  */
  assign n2462 = x_d1 == 9'b001010100;
  /* fplog32.vhdl:1335:50  */
  assign n2465 = x_d1 == 9'b001010101;
  /* fplog32.vhdl:1336:50  */
  assign n2468 = x_d1 == 9'b001010110;
  /* fplog32.vhdl:1337:50  */
  assign n2471 = x_d1 == 9'b001010111;
  /* fplog32.vhdl:1338:50  */
  assign n2474 = x_d1 == 9'b001011000;
  /* fplog32.vhdl:1339:50  */
  assign n2477 = x_d1 == 9'b001011001;
  /* fplog32.vhdl:1340:50  */
  assign n2480 = x_d1 == 9'b001011010;
  /* fplog32.vhdl:1341:50  */
  assign n2483 = x_d1 == 9'b001011011;
  /* fplog32.vhdl:1342:50  */
  assign n2486 = x_d1 == 9'b001011100;
  /* fplog32.vhdl:1343:50  */
  assign n2489 = x_d1 == 9'b001011101;
  /* fplog32.vhdl:1344:50  */
  assign n2492 = x_d1 == 9'b001011110;
  /* fplog32.vhdl:1345:50  */
  assign n2495 = x_d1 == 9'b001011111;
  /* fplog32.vhdl:1346:50  */
  assign n2498 = x_d1 == 9'b001100000;
  /* fplog32.vhdl:1347:50  */
  assign n2501 = x_d1 == 9'b001100001;
  /* fplog32.vhdl:1348:50  */
  assign n2504 = x_d1 == 9'b001100010;
  /* fplog32.vhdl:1349:50  */
  assign n2507 = x_d1 == 9'b001100011;
  /* fplog32.vhdl:1350:50  */
  assign n2510 = x_d1 == 9'b001100100;
  /* fplog32.vhdl:1351:50  */
  assign n2513 = x_d1 == 9'b001100101;
  /* fplog32.vhdl:1352:50  */
  assign n2516 = x_d1 == 9'b001100110;
  /* fplog32.vhdl:1353:50  */
  assign n2519 = x_d1 == 9'b001100111;
  /* fplog32.vhdl:1354:50  */
  assign n2522 = x_d1 == 9'b001101000;
  /* fplog32.vhdl:1355:50  */
  assign n2525 = x_d1 == 9'b001101001;
  /* fplog32.vhdl:1356:50  */
  assign n2528 = x_d1 == 9'b001101010;
  /* fplog32.vhdl:1357:50  */
  assign n2531 = x_d1 == 9'b001101011;
  /* fplog32.vhdl:1358:50  */
  assign n2534 = x_d1 == 9'b001101100;
  /* fplog32.vhdl:1359:50  */
  assign n2537 = x_d1 == 9'b001101101;
  /* fplog32.vhdl:1360:50  */
  assign n2540 = x_d1 == 9'b001101110;
  /* fplog32.vhdl:1361:50  */
  assign n2543 = x_d1 == 9'b001101111;
  /* fplog32.vhdl:1362:50  */
  assign n2546 = x_d1 == 9'b001110000;
  /* fplog32.vhdl:1363:50  */
  assign n2549 = x_d1 == 9'b001110001;
  /* fplog32.vhdl:1364:50  */
  assign n2552 = x_d1 == 9'b001110010;
  /* fplog32.vhdl:1365:50  */
  assign n2555 = x_d1 == 9'b001110011;
  /* fplog32.vhdl:1366:50  */
  assign n2558 = x_d1 == 9'b001110100;
  /* fplog32.vhdl:1367:50  */
  assign n2561 = x_d1 == 9'b001110101;
  /* fplog32.vhdl:1368:50  */
  assign n2564 = x_d1 == 9'b001110110;
  /* fplog32.vhdl:1369:50  */
  assign n2567 = x_d1 == 9'b001110111;
  /* fplog32.vhdl:1370:50  */
  assign n2570 = x_d1 == 9'b001111000;
  /* fplog32.vhdl:1371:50  */
  assign n2573 = x_d1 == 9'b001111001;
  /* fplog32.vhdl:1372:50  */
  assign n2576 = x_d1 == 9'b001111010;
  /* fplog32.vhdl:1373:50  */
  assign n2579 = x_d1 == 9'b001111011;
  /* fplog32.vhdl:1374:50  */
  assign n2582 = x_d1 == 9'b001111100;
  /* fplog32.vhdl:1375:50  */
  assign n2585 = x_d1 == 9'b001111101;
  /* fplog32.vhdl:1376:50  */
  assign n2588 = x_d1 == 9'b001111110;
  /* fplog32.vhdl:1377:50  */
  assign n2591 = x_d1 == 9'b001111111;
  /* fplog32.vhdl:1378:50  */
  assign n2594 = x_d1 == 9'b010000000;
  /* fplog32.vhdl:1379:50  */
  assign n2597 = x_d1 == 9'b010000001;
  /* fplog32.vhdl:1380:50  */
  assign n2600 = x_d1 == 9'b010000010;
  /* fplog32.vhdl:1381:50  */
  assign n2603 = x_d1 == 9'b010000011;
  /* fplog32.vhdl:1382:50  */
  assign n2606 = x_d1 == 9'b010000100;
  /* fplog32.vhdl:1383:50  */
  assign n2609 = x_d1 == 9'b010000101;
  /* fplog32.vhdl:1384:50  */
  assign n2612 = x_d1 == 9'b010000110;
  /* fplog32.vhdl:1385:50  */
  assign n2615 = x_d1 == 9'b010000111;
  /* fplog32.vhdl:1386:50  */
  assign n2618 = x_d1 == 9'b010001000;
  /* fplog32.vhdl:1387:50  */
  assign n2621 = x_d1 == 9'b010001001;
  /* fplog32.vhdl:1388:50  */
  assign n2624 = x_d1 == 9'b010001010;
  /* fplog32.vhdl:1389:50  */
  assign n2627 = x_d1 == 9'b010001011;
  /* fplog32.vhdl:1390:50  */
  assign n2630 = x_d1 == 9'b010001100;
  /* fplog32.vhdl:1391:50  */
  assign n2633 = x_d1 == 9'b010001101;
  /* fplog32.vhdl:1392:50  */
  assign n2636 = x_d1 == 9'b010001110;
  /* fplog32.vhdl:1393:50  */
  assign n2639 = x_d1 == 9'b010001111;
  /* fplog32.vhdl:1394:50  */
  assign n2642 = x_d1 == 9'b010010000;
  /* fplog32.vhdl:1395:50  */
  assign n2645 = x_d1 == 9'b010010001;
  /* fplog32.vhdl:1396:50  */
  assign n2648 = x_d1 == 9'b010010010;
  /* fplog32.vhdl:1397:50  */
  assign n2651 = x_d1 == 9'b010010011;
  /* fplog32.vhdl:1398:50  */
  assign n2654 = x_d1 == 9'b010010100;
  /* fplog32.vhdl:1399:50  */
  assign n2657 = x_d1 == 9'b010010101;
  /* fplog32.vhdl:1400:50  */
  assign n2660 = x_d1 == 9'b010010110;
  /* fplog32.vhdl:1401:50  */
  assign n2663 = x_d1 == 9'b010010111;
  /* fplog32.vhdl:1402:50  */
  assign n2666 = x_d1 == 9'b010011000;
  /* fplog32.vhdl:1403:50  */
  assign n2669 = x_d1 == 9'b010011001;
  /* fplog32.vhdl:1404:50  */
  assign n2672 = x_d1 == 9'b010011010;
  /* fplog32.vhdl:1405:50  */
  assign n2675 = x_d1 == 9'b010011011;
  /* fplog32.vhdl:1406:50  */
  assign n2678 = x_d1 == 9'b010011100;
  /* fplog32.vhdl:1407:50  */
  assign n2681 = x_d1 == 9'b010011101;
  /* fplog32.vhdl:1408:50  */
  assign n2684 = x_d1 == 9'b010011110;
  /* fplog32.vhdl:1409:50  */
  assign n2687 = x_d1 == 9'b010011111;
  /* fplog32.vhdl:1410:50  */
  assign n2690 = x_d1 == 9'b010100000;
  /* fplog32.vhdl:1411:50  */
  assign n2693 = x_d1 == 9'b010100001;
  /* fplog32.vhdl:1412:50  */
  assign n2696 = x_d1 == 9'b010100010;
  /* fplog32.vhdl:1413:50  */
  assign n2699 = x_d1 == 9'b010100011;
  /* fplog32.vhdl:1414:50  */
  assign n2702 = x_d1 == 9'b010100100;
  /* fplog32.vhdl:1415:50  */
  assign n2705 = x_d1 == 9'b010100101;
  /* fplog32.vhdl:1416:50  */
  assign n2708 = x_d1 == 9'b010100110;
  /* fplog32.vhdl:1417:50  */
  assign n2711 = x_d1 == 9'b010100111;
  /* fplog32.vhdl:1418:50  */
  assign n2714 = x_d1 == 9'b010101000;
  /* fplog32.vhdl:1419:50  */
  assign n2717 = x_d1 == 9'b010101001;
  /* fplog32.vhdl:1420:50  */
  assign n2720 = x_d1 == 9'b010101010;
  /* fplog32.vhdl:1421:50  */
  assign n2723 = x_d1 == 9'b010101011;
  /* fplog32.vhdl:1422:50  */
  assign n2726 = x_d1 == 9'b010101100;
  /* fplog32.vhdl:1423:50  */
  assign n2729 = x_d1 == 9'b010101101;
  /* fplog32.vhdl:1424:50  */
  assign n2732 = x_d1 == 9'b010101110;
  /* fplog32.vhdl:1425:50  */
  assign n2735 = x_d1 == 9'b010101111;
  /* fplog32.vhdl:1426:50  */
  assign n2738 = x_d1 == 9'b010110000;
  /* fplog32.vhdl:1427:50  */
  assign n2741 = x_d1 == 9'b010110001;
  /* fplog32.vhdl:1428:50  */
  assign n2744 = x_d1 == 9'b010110010;
  /* fplog32.vhdl:1429:50  */
  assign n2747 = x_d1 == 9'b010110011;
  /* fplog32.vhdl:1430:50  */
  assign n2750 = x_d1 == 9'b010110100;
  /* fplog32.vhdl:1431:50  */
  assign n2753 = x_d1 == 9'b010110101;
  /* fplog32.vhdl:1432:50  */
  assign n2756 = x_d1 == 9'b010110110;
  /* fplog32.vhdl:1433:50  */
  assign n2759 = x_d1 == 9'b010110111;
  /* fplog32.vhdl:1434:50  */
  assign n2762 = x_d1 == 9'b010111000;
  /* fplog32.vhdl:1435:50  */
  assign n2765 = x_d1 == 9'b010111001;
  /* fplog32.vhdl:1436:50  */
  assign n2768 = x_d1 == 9'b010111010;
  /* fplog32.vhdl:1437:50  */
  assign n2771 = x_d1 == 9'b010111011;
  /* fplog32.vhdl:1438:50  */
  assign n2774 = x_d1 == 9'b010111100;
  /* fplog32.vhdl:1439:50  */
  assign n2777 = x_d1 == 9'b010111101;
  /* fplog32.vhdl:1440:50  */
  assign n2780 = x_d1 == 9'b010111110;
  /* fplog32.vhdl:1441:50  */
  assign n2783 = x_d1 == 9'b010111111;
  /* fplog32.vhdl:1442:50  */
  assign n2786 = x_d1 == 9'b011000000;
  /* fplog32.vhdl:1443:50  */
  assign n2789 = x_d1 == 9'b011000001;
  /* fplog32.vhdl:1444:50  */
  assign n2792 = x_d1 == 9'b011000010;
  /* fplog32.vhdl:1445:50  */
  assign n2795 = x_d1 == 9'b011000011;
  /* fplog32.vhdl:1446:50  */
  assign n2798 = x_d1 == 9'b011000100;
  /* fplog32.vhdl:1447:50  */
  assign n2801 = x_d1 == 9'b011000101;
  /* fplog32.vhdl:1448:50  */
  assign n2804 = x_d1 == 9'b011000110;
  /* fplog32.vhdl:1449:50  */
  assign n2807 = x_d1 == 9'b011000111;
  /* fplog32.vhdl:1450:50  */
  assign n2810 = x_d1 == 9'b011001000;
  /* fplog32.vhdl:1451:50  */
  assign n2813 = x_d1 == 9'b011001001;
  /* fplog32.vhdl:1452:50  */
  assign n2816 = x_d1 == 9'b011001010;
  /* fplog32.vhdl:1453:50  */
  assign n2819 = x_d1 == 9'b011001011;
  /* fplog32.vhdl:1454:50  */
  assign n2822 = x_d1 == 9'b011001100;
  /* fplog32.vhdl:1455:50  */
  assign n2825 = x_d1 == 9'b011001101;
  /* fplog32.vhdl:1456:50  */
  assign n2828 = x_d1 == 9'b011001110;
  /* fplog32.vhdl:1457:50  */
  assign n2831 = x_d1 == 9'b011001111;
  /* fplog32.vhdl:1458:50  */
  assign n2834 = x_d1 == 9'b011010000;
  /* fplog32.vhdl:1459:50  */
  assign n2837 = x_d1 == 9'b011010001;
  /* fplog32.vhdl:1460:50  */
  assign n2840 = x_d1 == 9'b011010010;
  /* fplog32.vhdl:1461:50  */
  assign n2843 = x_d1 == 9'b011010011;
  /* fplog32.vhdl:1462:50  */
  assign n2846 = x_d1 == 9'b011010100;
  /* fplog32.vhdl:1463:50  */
  assign n2849 = x_d1 == 9'b011010101;
  /* fplog32.vhdl:1464:50  */
  assign n2852 = x_d1 == 9'b011010110;
  /* fplog32.vhdl:1465:50  */
  assign n2855 = x_d1 == 9'b011010111;
  /* fplog32.vhdl:1466:50  */
  assign n2858 = x_d1 == 9'b011011000;
  /* fplog32.vhdl:1467:50  */
  assign n2861 = x_d1 == 9'b011011001;
  /* fplog32.vhdl:1468:50  */
  assign n2864 = x_d1 == 9'b011011010;
  /* fplog32.vhdl:1469:50  */
  assign n2867 = x_d1 == 9'b011011011;
  /* fplog32.vhdl:1470:50  */
  assign n2870 = x_d1 == 9'b011011100;
  /* fplog32.vhdl:1471:50  */
  assign n2873 = x_d1 == 9'b011011101;
  /* fplog32.vhdl:1472:50  */
  assign n2876 = x_d1 == 9'b011011110;
  /* fplog32.vhdl:1473:50  */
  assign n2879 = x_d1 == 9'b011011111;
  /* fplog32.vhdl:1474:50  */
  assign n2882 = x_d1 == 9'b011100000;
  /* fplog32.vhdl:1475:50  */
  assign n2885 = x_d1 == 9'b011100001;
  /* fplog32.vhdl:1476:50  */
  assign n2888 = x_d1 == 9'b011100010;
  /* fplog32.vhdl:1477:50  */
  assign n2891 = x_d1 == 9'b011100011;
  /* fplog32.vhdl:1478:50  */
  assign n2894 = x_d1 == 9'b011100100;
  /* fplog32.vhdl:1479:50  */
  assign n2897 = x_d1 == 9'b011100101;
  /* fplog32.vhdl:1480:50  */
  assign n2900 = x_d1 == 9'b011100110;
  /* fplog32.vhdl:1481:50  */
  assign n2903 = x_d1 == 9'b011100111;
  /* fplog32.vhdl:1482:50  */
  assign n2906 = x_d1 == 9'b011101000;
  /* fplog32.vhdl:1483:50  */
  assign n2909 = x_d1 == 9'b011101001;
  /* fplog32.vhdl:1484:50  */
  assign n2912 = x_d1 == 9'b011101010;
  /* fplog32.vhdl:1485:50  */
  assign n2915 = x_d1 == 9'b011101011;
  /* fplog32.vhdl:1486:50  */
  assign n2918 = x_d1 == 9'b011101100;
  /* fplog32.vhdl:1487:50  */
  assign n2921 = x_d1 == 9'b011101101;
  /* fplog32.vhdl:1488:50  */
  assign n2924 = x_d1 == 9'b011101110;
  /* fplog32.vhdl:1489:50  */
  assign n2927 = x_d1 == 9'b011101111;
  /* fplog32.vhdl:1490:50  */
  assign n2930 = x_d1 == 9'b011110000;
  /* fplog32.vhdl:1491:50  */
  assign n2933 = x_d1 == 9'b011110001;
  /* fplog32.vhdl:1492:50  */
  assign n2936 = x_d1 == 9'b011110010;
  /* fplog32.vhdl:1493:50  */
  assign n2939 = x_d1 == 9'b011110011;
  /* fplog32.vhdl:1494:50  */
  assign n2942 = x_d1 == 9'b011110100;
  /* fplog32.vhdl:1495:50  */
  assign n2945 = x_d1 == 9'b011110101;
  /* fplog32.vhdl:1496:50  */
  assign n2948 = x_d1 == 9'b011110110;
  /* fplog32.vhdl:1497:50  */
  assign n2951 = x_d1 == 9'b011110111;
  /* fplog32.vhdl:1498:50  */
  assign n2954 = x_d1 == 9'b011111000;
  /* fplog32.vhdl:1499:50  */
  assign n2957 = x_d1 == 9'b011111001;
  /* fplog32.vhdl:1500:50  */
  assign n2960 = x_d1 == 9'b011111010;
  /* fplog32.vhdl:1501:50  */
  assign n2963 = x_d1 == 9'b011111011;
  /* fplog32.vhdl:1502:50  */
  assign n2966 = x_d1 == 9'b011111100;
  /* fplog32.vhdl:1503:50  */
  assign n2969 = x_d1 == 9'b011111101;
  /* fplog32.vhdl:1504:50  */
  assign n2972 = x_d1 == 9'b011111110;
  /* fplog32.vhdl:1505:50  */
  assign n2975 = x_d1 == 9'b011111111;
  /* fplog32.vhdl:1506:50  */
  assign n2978 = x_d1 == 9'b100000000;
  /* fplog32.vhdl:1507:50  */
  assign n2981 = x_d1 == 9'b100000001;
  /* fplog32.vhdl:1508:50  */
  assign n2984 = x_d1 == 9'b100000010;
  /* fplog32.vhdl:1509:50  */
  assign n2987 = x_d1 == 9'b100000011;
  /* fplog32.vhdl:1510:50  */
  assign n2990 = x_d1 == 9'b100000100;
  /* fplog32.vhdl:1511:50  */
  assign n2993 = x_d1 == 9'b100000101;
  /* fplog32.vhdl:1512:50  */
  assign n2996 = x_d1 == 9'b100000110;
  /* fplog32.vhdl:1513:50  */
  assign n2999 = x_d1 == 9'b100000111;
  /* fplog32.vhdl:1514:50  */
  assign n3002 = x_d1 == 9'b100001000;
  /* fplog32.vhdl:1515:50  */
  assign n3005 = x_d1 == 9'b100001001;
  /* fplog32.vhdl:1516:50  */
  assign n3008 = x_d1 == 9'b100001010;
  /* fplog32.vhdl:1517:50  */
  assign n3011 = x_d1 == 9'b100001011;
  /* fplog32.vhdl:1518:50  */
  assign n3014 = x_d1 == 9'b100001100;
  /* fplog32.vhdl:1519:50  */
  assign n3017 = x_d1 == 9'b100001101;
  /* fplog32.vhdl:1520:50  */
  assign n3020 = x_d1 == 9'b100001110;
  /* fplog32.vhdl:1521:50  */
  assign n3023 = x_d1 == 9'b100001111;
  /* fplog32.vhdl:1522:50  */
  assign n3026 = x_d1 == 9'b100010000;
  /* fplog32.vhdl:1523:50  */
  assign n3029 = x_d1 == 9'b100010001;
  /* fplog32.vhdl:1524:50  */
  assign n3032 = x_d1 == 9'b100010010;
  /* fplog32.vhdl:1525:50  */
  assign n3035 = x_d1 == 9'b100010011;
  /* fplog32.vhdl:1526:50  */
  assign n3038 = x_d1 == 9'b100010100;
  /* fplog32.vhdl:1527:50  */
  assign n3041 = x_d1 == 9'b100010101;
  /* fplog32.vhdl:1528:50  */
  assign n3044 = x_d1 == 9'b100010110;
  /* fplog32.vhdl:1529:50  */
  assign n3047 = x_d1 == 9'b100010111;
  /* fplog32.vhdl:1530:50  */
  assign n3050 = x_d1 == 9'b100011000;
  /* fplog32.vhdl:1531:50  */
  assign n3053 = x_d1 == 9'b100011001;
  /* fplog32.vhdl:1532:50  */
  assign n3056 = x_d1 == 9'b100011010;
  /* fplog32.vhdl:1533:50  */
  assign n3059 = x_d1 == 9'b100011011;
  /* fplog32.vhdl:1534:50  */
  assign n3062 = x_d1 == 9'b100011100;
  /* fplog32.vhdl:1535:50  */
  assign n3065 = x_d1 == 9'b100011101;
  /* fplog32.vhdl:1536:50  */
  assign n3068 = x_d1 == 9'b100011110;
  /* fplog32.vhdl:1537:50  */
  assign n3071 = x_d1 == 9'b100011111;
  /* fplog32.vhdl:1538:50  */
  assign n3074 = x_d1 == 9'b100100000;
  /* fplog32.vhdl:1539:50  */
  assign n3077 = x_d1 == 9'b100100001;
  /* fplog32.vhdl:1540:50  */
  assign n3080 = x_d1 == 9'b100100010;
  /* fplog32.vhdl:1541:50  */
  assign n3083 = x_d1 == 9'b100100011;
  /* fplog32.vhdl:1542:50  */
  assign n3086 = x_d1 == 9'b100100100;
  /* fplog32.vhdl:1543:50  */
  assign n3089 = x_d1 == 9'b100100101;
  /* fplog32.vhdl:1544:50  */
  assign n3092 = x_d1 == 9'b100100110;
  /* fplog32.vhdl:1545:50  */
  assign n3095 = x_d1 == 9'b100100111;
  /* fplog32.vhdl:1546:50  */
  assign n3098 = x_d1 == 9'b100101000;
  /* fplog32.vhdl:1547:50  */
  assign n3101 = x_d1 == 9'b100101001;
  /* fplog32.vhdl:1548:50  */
  assign n3104 = x_d1 == 9'b100101010;
  /* fplog32.vhdl:1549:50  */
  assign n3107 = x_d1 == 9'b100101011;
  /* fplog32.vhdl:1550:50  */
  assign n3110 = x_d1 == 9'b100101100;
  /* fplog32.vhdl:1551:50  */
  assign n3113 = x_d1 == 9'b100101101;
  /* fplog32.vhdl:1552:50  */
  assign n3116 = x_d1 == 9'b100101110;
  /* fplog32.vhdl:1553:50  */
  assign n3119 = x_d1 == 9'b100101111;
  /* fplog32.vhdl:1554:50  */
  assign n3122 = x_d1 == 9'b100110000;
  /* fplog32.vhdl:1555:50  */
  assign n3125 = x_d1 == 9'b100110001;
  /* fplog32.vhdl:1556:50  */
  assign n3128 = x_d1 == 9'b100110010;
  /* fplog32.vhdl:1557:50  */
  assign n3131 = x_d1 == 9'b100110011;
  /* fplog32.vhdl:1558:50  */
  assign n3134 = x_d1 == 9'b100110100;
  /* fplog32.vhdl:1559:50  */
  assign n3137 = x_d1 == 9'b100110101;
  /* fplog32.vhdl:1560:50  */
  assign n3140 = x_d1 == 9'b100110110;
  /* fplog32.vhdl:1561:50  */
  assign n3143 = x_d1 == 9'b100110111;
  /* fplog32.vhdl:1562:50  */
  assign n3146 = x_d1 == 9'b100111000;
  /* fplog32.vhdl:1563:50  */
  assign n3149 = x_d1 == 9'b100111001;
  /* fplog32.vhdl:1564:50  */
  assign n3152 = x_d1 == 9'b100111010;
  /* fplog32.vhdl:1565:50  */
  assign n3155 = x_d1 == 9'b100111011;
  /* fplog32.vhdl:1566:50  */
  assign n3158 = x_d1 == 9'b100111100;
  /* fplog32.vhdl:1567:50  */
  assign n3161 = x_d1 == 9'b100111101;
  /* fplog32.vhdl:1568:50  */
  assign n3164 = x_d1 == 9'b100111110;
  /* fplog32.vhdl:1569:50  */
  assign n3167 = x_d1 == 9'b100111111;
  /* fplog32.vhdl:1570:50  */
  assign n3170 = x_d1 == 9'b101000000;
  /* fplog32.vhdl:1571:50  */
  assign n3173 = x_d1 == 9'b101000001;
  /* fplog32.vhdl:1572:50  */
  assign n3176 = x_d1 == 9'b101000010;
  /* fplog32.vhdl:1573:50  */
  assign n3179 = x_d1 == 9'b101000011;
  /* fplog32.vhdl:1574:50  */
  assign n3182 = x_d1 == 9'b101000100;
  /* fplog32.vhdl:1575:50  */
  assign n3185 = x_d1 == 9'b101000101;
  /* fplog32.vhdl:1576:50  */
  assign n3188 = x_d1 == 9'b101000110;
  /* fplog32.vhdl:1577:50  */
  assign n3191 = x_d1 == 9'b101000111;
  /* fplog32.vhdl:1578:50  */
  assign n3194 = x_d1 == 9'b101001000;
  /* fplog32.vhdl:1579:50  */
  assign n3197 = x_d1 == 9'b101001001;
  /* fplog32.vhdl:1580:50  */
  assign n3200 = x_d1 == 9'b101001010;
  /* fplog32.vhdl:1581:50  */
  assign n3203 = x_d1 == 9'b101001011;
  /* fplog32.vhdl:1582:50  */
  assign n3206 = x_d1 == 9'b101001100;
  /* fplog32.vhdl:1583:50  */
  assign n3209 = x_d1 == 9'b101001101;
  /* fplog32.vhdl:1584:50  */
  assign n3212 = x_d1 == 9'b101001110;
  /* fplog32.vhdl:1585:50  */
  assign n3215 = x_d1 == 9'b101001111;
  /* fplog32.vhdl:1586:50  */
  assign n3218 = x_d1 == 9'b101010000;
  /* fplog32.vhdl:1587:50  */
  assign n3221 = x_d1 == 9'b101010001;
  /* fplog32.vhdl:1588:50  */
  assign n3224 = x_d1 == 9'b101010010;
  /* fplog32.vhdl:1589:50  */
  assign n3227 = x_d1 == 9'b101010011;
  /* fplog32.vhdl:1590:50  */
  assign n3230 = x_d1 == 9'b101010100;
  /* fplog32.vhdl:1591:50  */
  assign n3233 = x_d1 == 9'b101010101;
  /* fplog32.vhdl:1592:50  */
  assign n3236 = x_d1 == 9'b101010110;
  /* fplog32.vhdl:1593:50  */
  assign n3239 = x_d1 == 9'b101010111;
  /* fplog32.vhdl:1594:50  */
  assign n3242 = x_d1 == 9'b101011000;
  /* fplog32.vhdl:1595:50  */
  assign n3245 = x_d1 == 9'b101011001;
  /* fplog32.vhdl:1596:50  */
  assign n3248 = x_d1 == 9'b101011010;
  /* fplog32.vhdl:1597:50  */
  assign n3251 = x_d1 == 9'b101011011;
  /* fplog32.vhdl:1598:50  */
  assign n3254 = x_d1 == 9'b101011100;
  /* fplog32.vhdl:1599:50  */
  assign n3257 = x_d1 == 9'b101011101;
  /* fplog32.vhdl:1600:50  */
  assign n3260 = x_d1 == 9'b101011110;
  /* fplog32.vhdl:1601:50  */
  assign n3263 = x_d1 == 9'b101011111;
  /* fplog32.vhdl:1602:50  */
  assign n3266 = x_d1 == 9'b101100000;
  /* fplog32.vhdl:1603:50  */
  assign n3269 = x_d1 == 9'b101100001;
  /* fplog32.vhdl:1604:50  */
  assign n3272 = x_d1 == 9'b101100010;
  /* fplog32.vhdl:1605:50  */
  assign n3275 = x_d1 == 9'b101100011;
  /* fplog32.vhdl:1606:50  */
  assign n3278 = x_d1 == 9'b101100100;
  /* fplog32.vhdl:1607:50  */
  assign n3281 = x_d1 == 9'b101100101;
  /* fplog32.vhdl:1608:50  */
  assign n3284 = x_d1 == 9'b101100110;
  /* fplog32.vhdl:1609:50  */
  assign n3287 = x_d1 == 9'b101100111;
  /* fplog32.vhdl:1610:50  */
  assign n3290 = x_d1 == 9'b101101000;
  /* fplog32.vhdl:1611:50  */
  assign n3293 = x_d1 == 9'b101101001;
  /* fplog32.vhdl:1612:50  */
  assign n3296 = x_d1 == 9'b101101010;
  /* fplog32.vhdl:1613:50  */
  assign n3299 = x_d1 == 9'b101101011;
  /* fplog32.vhdl:1614:50  */
  assign n3302 = x_d1 == 9'b101101100;
  /* fplog32.vhdl:1615:50  */
  assign n3305 = x_d1 == 9'b101101101;
  /* fplog32.vhdl:1616:50  */
  assign n3308 = x_d1 == 9'b101101110;
  /* fplog32.vhdl:1617:50  */
  assign n3311 = x_d1 == 9'b101101111;
  /* fplog32.vhdl:1618:50  */
  assign n3314 = x_d1 == 9'b101110000;
  /* fplog32.vhdl:1619:50  */
  assign n3317 = x_d1 == 9'b101110001;
  /* fplog32.vhdl:1620:50  */
  assign n3320 = x_d1 == 9'b101110010;
  /* fplog32.vhdl:1621:50  */
  assign n3323 = x_d1 == 9'b101110011;
  /* fplog32.vhdl:1622:50  */
  assign n3326 = x_d1 == 9'b101110100;
  /* fplog32.vhdl:1623:50  */
  assign n3329 = x_d1 == 9'b101110101;
  /* fplog32.vhdl:1624:50  */
  assign n3332 = x_d1 == 9'b101110110;
  /* fplog32.vhdl:1625:50  */
  assign n3335 = x_d1 == 9'b101110111;
  /* fplog32.vhdl:1626:50  */
  assign n3338 = x_d1 == 9'b101111000;
  /* fplog32.vhdl:1627:50  */
  assign n3341 = x_d1 == 9'b101111001;
  /* fplog32.vhdl:1628:50  */
  assign n3344 = x_d1 == 9'b101111010;
  /* fplog32.vhdl:1629:50  */
  assign n3347 = x_d1 == 9'b101111011;
  /* fplog32.vhdl:1630:50  */
  assign n3350 = x_d1 == 9'b101111100;
  /* fplog32.vhdl:1631:50  */
  assign n3353 = x_d1 == 9'b101111101;
  /* fplog32.vhdl:1632:50  */
  assign n3356 = x_d1 == 9'b101111110;
  /* fplog32.vhdl:1633:50  */
  assign n3359 = x_d1 == 9'b101111111;
  /* fplog32.vhdl:1634:50  */
  assign n3362 = x_d1 == 9'b110000000;
  /* fplog32.vhdl:1635:50  */
  assign n3365 = x_d1 == 9'b110000001;
  /* fplog32.vhdl:1636:50  */
  assign n3368 = x_d1 == 9'b110000010;
  /* fplog32.vhdl:1637:50  */
  assign n3371 = x_d1 == 9'b110000011;
  /* fplog32.vhdl:1638:50  */
  assign n3374 = x_d1 == 9'b110000100;
  /* fplog32.vhdl:1639:50  */
  assign n3377 = x_d1 == 9'b110000101;
  /* fplog32.vhdl:1640:50  */
  assign n3380 = x_d1 == 9'b110000110;
  /* fplog32.vhdl:1641:50  */
  assign n3383 = x_d1 == 9'b110000111;
  /* fplog32.vhdl:1642:50  */
  assign n3386 = x_d1 == 9'b110001000;
  /* fplog32.vhdl:1643:50  */
  assign n3389 = x_d1 == 9'b110001001;
  /* fplog32.vhdl:1644:50  */
  assign n3392 = x_d1 == 9'b110001010;
  /* fplog32.vhdl:1645:50  */
  assign n3395 = x_d1 == 9'b110001011;
  /* fplog32.vhdl:1646:50  */
  assign n3398 = x_d1 == 9'b110001100;
  /* fplog32.vhdl:1647:50  */
  assign n3401 = x_d1 == 9'b110001101;
  /* fplog32.vhdl:1648:50  */
  assign n3404 = x_d1 == 9'b110001110;
  /* fplog32.vhdl:1649:50  */
  assign n3407 = x_d1 == 9'b110001111;
  /* fplog32.vhdl:1650:50  */
  assign n3410 = x_d1 == 9'b110010000;
  /* fplog32.vhdl:1651:50  */
  assign n3413 = x_d1 == 9'b110010001;
  /* fplog32.vhdl:1652:50  */
  assign n3416 = x_d1 == 9'b110010010;
  /* fplog32.vhdl:1653:50  */
  assign n3419 = x_d1 == 9'b110010011;
  /* fplog32.vhdl:1654:50  */
  assign n3422 = x_d1 == 9'b110010100;
  /* fplog32.vhdl:1655:50  */
  assign n3425 = x_d1 == 9'b110010101;
  /* fplog32.vhdl:1656:50  */
  assign n3428 = x_d1 == 9'b110010110;
  /* fplog32.vhdl:1657:50  */
  assign n3431 = x_d1 == 9'b110010111;
  /* fplog32.vhdl:1658:50  */
  assign n3434 = x_d1 == 9'b110011000;
  /* fplog32.vhdl:1659:50  */
  assign n3437 = x_d1 == 9'b110011001;
  /* fplog32.vhdl:1660:50  */
  assign n3440 = x_d1 == 9'b110011010;
  /* fplog32.vhdl:1661:50  */
  assign n3443 = x_d1 == 9'b110011011;
  /* fplog32.vhdl:1662:50  */
  assign n3446 = x_d1 == 9'b110011100;
  /* fplog32.vhdl:1663:50  */
  assign n3449 = x_d1 == 9'b110011101;
  /* fplog32.vhdl:1664:50  */
  assign n3452 = x_d1 == 9'b110011110;
  /* fplog32.vhdl:1665:50  */
  assign n3455 = x_d1 == 9'b110011111;
  /* fplog32.vhdl:1666:50  */
  assign n3458 = x_d1 == 9'b110100000;
  /* fplog32.vhdl:1667:50  */
  assign n3461 = x_d1 == 9'b110100001;
  /* fplog32.vhdl:1668:50  */
  assign n3464 = x_d1 == 9'b110100010;
  /* fplog32.vhdl:1669:50  */
  assign n3467 = x_d1 == 9'b110100011;
  /* fplog32.vhdl:1670:50  */
  assign n3470 = x_d1 == 9'b110100100;
  /* fplog32.vhdl:1671:50  */
  assign n3473 = x_d1 == 9'b110100101;
  /* fplog32.vhdl:1672:50  */
  assign n3476 = x_d1 == 9'b110100110;
  /* fplog32.vhdl:1673:50  */
  assign n3479 = x_d1 == 9'b110100111;
  /* fplog32.vhdl:1674:50  */
  assign n3482 = x_d1 == 9'b110101000;
  /* fplog32.vhdl:1675:50  */
  assign n3485 = x_d1 == 9'b110101001;
  /* fplog32.vhdl:1676:50  */
  assign n3488 = x_d1 == 9'b110101010;
  /* fplog32.vhdl:1677:50  */
  assign n3491 = x_d1 == 9'b110101011;
  /* fplog32.vhdl:1678:50  */
  assign n3494 = x_d1 == 9'b110101100;
  /* fplog32.vhdl:1679:50  */
  assign n3497 = x_d1 == 9'b110101101;
  /* fplog32.vhdl:1680:50  */
  assign n3500 = x_d1 == 9'b110101110;
  /* fplog32.vhdl:1681:50  */
  assign n3503 = x_d1 == 9'b110101111;
  /* fplog32.vhdl:1682:50  */
  assign n3506 = x_d1 == 9'b110110000;
  /* fplog32.vhdl:1683:50  */
  assign n3509 = x_d1 == 9'b110110001;
  /* fplog32.vhdl:1684:50  */
  assign n3512 = x_d1 == 9'b110110010;
  /* fplog32.vhdl:1685:50  */
  assign n3515 = x_d1 == 9'b110110011;
  /* fplog32.vhdl:1686:50  */
  assign n3518 = x_d1 == 9'b110110100;
  /* fplog32.vhdl:1687:50  */
  assign n3521 = x_d1 == 9'b110110101;
  /* fplog32.vhdl:1688:50  */
  assign n3524 = x_d1 == 9'b110110110;
  /* fplog32.vhdl:1689:50  */
  assign n3527 = x_d1 == 9'b110110111;
  /* fplog32.vhdl:1690:50  */
  assign n3530 = x_d1 == 9'b110111000;
  /* fplog32.vhdl:1691:50  */
  assign n3533 = x_d1 == 9'b110111001;
  /* fplog32.vhdl:1692:50  */
  assign n3536 = x_d1 == 9'b110111010;
  /* fplog32.vhdl:1693:50  */
  assign n3539 = x_d1 == 9'b110111011;
  /* fplog32.vhdl:1694:50  */
  assign n3542 = x_d1 == 9'b110111100;
  /* fplog32.vhdl:1695:50  */
  assign n3545 = x_d1 == 9'b110111101;
  /* fplog32.vhdl:1696:50  */
  assign n3548 = x_d1 == 9'b110111110;
  /* fplog32.vhdl:1697:50  */
  assign n3551 = x_d1 == 9'b110111111;
  /* fplog32.vhdl:1698:50  */
  assign n3554 = x_d1 == 9'b111000000;
  /* fplog32.vhdl:1699:50  */
  assign n3557 = x_d1 == 9'b111000001;
  /* fplog32.vhdl:1700:50  */
  assign n3560 = x_d1 == 9'b111000010;
  /* fplog32.vhdl:1701:50  */
  assign n3563 = x_d1 == 9'b111000011;
  /* fplog32.vhdl:1702:50  */
  assign n3566 = x_d1 == 9'b111000100;
  /* fplog32.vhdl:1703:50  */
  assign n3569 = x_d1 == 9'b111000101;
  /* fplog32.vhdl:1704:50  */
  assign n3572 = x_d1 == 9'b111000110;
  /* fplog32.vhdl:1705:50  */
  assign n3575 = x_d1 == 9'b111000111;
  /* fplog32.vhdl:1706:50  */
  assign n3578 = x_d1 == 9'b111001000;
  /* fplog32.vhdl:1707:50  */
  assign n3581 = x_d1 == 9'b111001001;
  /* fplog32.vhdl:1708:50  */
  assign n3584 = x_d1 == 9'b111001010;
  /* fplog32.vhdl:1709:50  */
  assign n3587 = x_d1 == 9'b111001011;
  /* fplog32.vhdl:1710:50  */
  assign n3590 = x_d1 == 9'b111001100;
  /* fplog32.vhdl:1711:50  */
  assign n3593 = x_d1 == 9'b111001101;
  /* fplog32.vhdl:1712:50  */
  assign n3596 = x_d1 == 9'b111001110;
  /* fplog32.vhdl:1713:50  */
  assign n3599 = x_d1 == 9'b111001111;
  /* fplog32.vhdl:1714:50  */
  assign n3602 = x_d1 == 9'b111010000;
  /* fplog32.vhdl:1715:50  */
  assign n3605 = x_d1 == 9'b111010001;
  /* fplog32.vhdl:1716:50  */
  assign n3608 = x_d1 == 9'b111010010;
  /* fplog32.vhdl:1717:50  */
  assign n3611 = x_d1 == 9'b111010011;
  /* fplog32.vhdl:1718:50  */
  assign n3614 = x_d1 == 9'b111010100;
  /* fplog32.vhdl:1719:50  */
  assign n3617 = x_d1 == 9'b111010101;
  /* fplog32.vhdl:1720:50  */
  assign n3620 = x_d1 == 9'b111010110;
  /* fplog32.vhdl:1721:50  */
  assign n3623 = x_d1 == 9'b111010111;
  /* fplog32.vhdl:1722:50  */
  assign n3626 = x_d1 == 9'b111011000;
  /* fplog32.vhdl:1723:50  */
  assign n3629 = x_d1 == 9'b111011001;
  /* fplog32.vhdl:1724:50  */
  assign n3632 = x_d1 == 9'b111011010;
  /* fplog32.vhdl:1725:50  */
  assign n3635 = x_d1 == 9'b111011011;
  /* fplog32.vhdl:1726:50  */
  assign n3638 = x_d1 == 9'b111011100;
  /* fplog32.vhdl:1727:50  */
  assign n3641 = x_d1 == 9'b111011101;
  /* fplog32.vhdl:1728:50  */
  assign n3644 = x_d1 == 9'b111011110;
  /* fplog32.vhdl:1729:50  */
  assign n3647 = x_d1 == 9'b111011111;
  /* fplog32.vhdl:1730:50  */
  assign n3650 = x_d1 == 9'b111100000;
  /* fplog32.vhdl:1731:50  */
  assign n3653 = x_d1 == 9'b111100001;
  /* fplog32.vhdl:1732:50  */
  assign n3656 = x_d1 == 9'b111100010;
  /* fplog32.vhdl:1733:50  */
  assign n3659 = x_d1 == 9'b111100011;
  /* fplog32.vhdl:1734:50  */
  assign n3662 = x_d1 == 9'b111100100;
  /* fplog32.vhdl:1735:50  */
  assign n3665 = x_d1 == 9'b111100101;
  /* fplog32.vhdl:1736:50  */
  assign n3668 = x_d1 == 9'b111100110;
  /* fplog32.vhdl:1737:50  */
  assign n3671 = x_d1 == 9'b111100111;
  /* fplog32.vhdl:1738:50  */
  assign n3674 = x_d1 == 9'b111101000;
  /* fplog32.vhdl:1739:50  */
  assign n3677 = x_d1 == 9'b111101001;
  /* fplog32.vhdl:1740:50  */
  assign n3680 = x_d1 == 9'b111101010;
  /* fplog32.vhdl:1741:50  */
  assign n3683 = x_d1 == 9'b111101011;
  /* fplog32.vhdl:1742:50  */
  assign n3686 = x_d1 == 9'b111101100;
  /* fplog32.vhdl:1743:50  */
  assign n3689 = x_d1 == 9'b111101101;
  /* fplog32.vhdl:1744:50  */
  assign n3692 = x_d1 == 9'b111101110;
  /* fplog32.vhdl:1745:50  */
  assign n3695 = x_d1 == 9'b111101111;
  /* fplog32.vhdl:1746:50  */
  assign n3698 = x_d1 == 9'b111110000;
  /* fplog32.vhdl:1747:50  */
  assign n3701 = x_d1 == 9'b111110001;
  /* fplog32.vhdl:1748:50  */
  assign n3704 = x_d1 == 9'b111110010;
  /* fplog32.vhdl:1749:50  */
  assign n3707 = x_d1 == 9'b111110011;
  /* fplog32.vhdl:1750:50  */
  assign n3710 = x_d1 == 9'b111110100;
  /* fplog32.vhdl:1751:50  */
  assign n3713 = x_d1 == 9'b111110101;
  /* fplog32.vhdl:1752:50  */
  assign n3716 = x_d1 == 9'b111110110;
  /* fplog32.vhdl:1753:50  */
  assign n3719 = x_d1 == 9'b111110111;
  /* fplog32.vhdl:1754:50  */
  assign n3722 = x_d1 == 9'b111111000;
  /* fplog32.vhdl:1755:50  */
  assign n3725 = x_d1 == 9'b111111001;
  /* fplog32.vhdl:1756:50  */
  assign n3728 = x_d1 == 9'b111111010;
  /* fplog32.vhdl:1757:50  */
  assign n3731 = x_d1 == 9'b111111011;
  /* fplog32.vhdl:1758:50  */
  assign n3734 = x_d1 == 9'b111111100;
  /* fplog32.vhdl:1759:50  */
  assign n3737 = x_d1 == 9'b111111101;
  /* fplog32.vhdl:1760:50  */
  assign n3740 = x_d1 == 9'b111111110;
  /* fplog32.vhdl:1761:50  */
  assign n3743 = x_d1 == 9'b111111111;
  assign n3745 = {n3743, n3740, n3737, n3734, n3731, n3728, n3725, n3722, n3719, n3716, n3713, n3710, n3707, n3704, n3701, n3698, n3695, n3692, n3689, n3686, n3683, n3680, n3677, n3674, n3671, n3668, n3665, n3662, n3659, n3656, n3653, n3650, n3647, n3644, n3641, n3638, n3635, n3632, n3629, n3626, n3623, n3620, n3617, n3614, n3611, n3608, n3605, n3602, n3599, n3596, n3593, n3590, n3587, n3584, n3581, n3578, n3575, n3572, n3569, n3566, n3563, n3560, n3557, n3554, n3551, n3548, n3545, n3542, n3539, n3536, n3533, n3530, n3527, n3524, n3521, n3518, n3515, n3512, n3509, n3506, n3503, n3500, n3497, n3494, n3491, n3488, n3485, n3482, n3479, n3476, n3473, n3470, n3467, n3464, n3461, n3458, n3455, n3452, n3449, n3446, n3443, n3440, n3437, n3434, n3431, n3428, n3425, n3422, n3419, n3416, n3413, n3410, n3407, n3404, n3401, n3398, n3395, n3392, n3389, n3386, n3383, n3380, n3377, n3374, n3371, n3368, n3365, n3362, n3359, n3356, n3353, n3350, n3347, n3344, n3341, n3338, n3335, n3332, n3329, n3326, n3323, n3320, n3317, n3314, n3311, n3308, n3305, n3302, n3299, n3296, n3293, n3290, n3287, n3284, n3281, n3278, n3275, n3272, n3269, n3266, n3263, n3260, n3257, n3254, n3251, n3248, n3245, n3242, n3239, n3236, n3233, n3230, n3227, n3224, n3221, n3218, n3215, n3212, n3209, n3206, n3203, n3200, n3197, n3194, n3191, n3188, n3185, n3182, n3179, n3176, n3173, n3170, n3167, n3164, n3161, n3158, n3155, n3152, n3149, n3146, n3143, n3140, n3137, n3134, n3131, n3128, n3125, n3122, n3119, n3116, n3113, n3110, n3107, n3104, n3101, n3098, n3095, n3092, n3089, n3086, n3083, n3080, n3077, n3074, n3071, n3068, n3065, n3062, n3059, n3056, n3053, n3050, n3047, n3044, n3041, n3038, n3035, n3032, n3029, n3026, n3023, n3020, n3017, n3014, n3011, n3008, n3005, n3002, n2999, n2996, n2993, n2990, n2987, n2984, n2981, n2978, n2975, n2972, n2969, n2966, n2963, n2960, n2957, n2954, n2951, n2948, n2945, n2942, n2939, n2936, n2933, n2930, n2927, n2924, n2921, n2918, n2915, n2912, n2909, n2906, n2903, n2900, n2897, n2894, n2891, n2888, n2885, n2882, n2879, n2876, n2873, n2870, n2867, n2864, n2861, n2858, n2855, n2852, n2849, n2846, n2843, n2840, n2837, n2834, n2831, n2828, n2825, n2822, n2819, n2816, n2813, n2810, n2807, n2804, n2801, n2798, n2795, n2792, n2789, n2786, n2783, n2780, n2777, n2774, n2771, n2768, n2765, n2762, n2759, n2756, n2753, n2750, n2747, n2744, n2741, n2738, n2735, n2732, n2729, n2726, n2723, n2720, n2717, n2714, n2711, n2708, n2705, n2702, n2699, n2696, n2693, n2690, n2687, n2684, n2681, n2678, n2675, n2672, n2669, n2666, n2663, n2660, n2657, n2654, n2651, n2648, n2645, n2642, n2639, n2636, n2633, n2630, n2627, n2624, n2621, n2618, n2615, n2612, n2609, n2606, n2603, n2600, n2597, n2594, n2591, n2588, n2585, n2582, n2579, n2576, n2573, n2570, n2567, n2564, n2561, n2558, n2555, n2552, n2549, n2546, n2543, n2540, n2537, n2534, n2531, n2528, n2525, n2522, n2519, n2516, n2513, n2510, n2507, n2504, n2501, n2498, n2495, n2492, n2489, n2486, n2483, n2480, n2477, n2474, n2471, n2468, n2465, n2462, n2459, n2456, n2453, n2450, n2447, n2444, n2441, n2438, n2435, n2432, n2429, n2426, n2423, n2420, n2417, n2414, n2411, n2408, n2405, n2402, n2399, n2396, n2393, n2390, n2387, n2384, n2381, n2378, n2375, n2372, n2369, n2366, n2363, n2360, n2357, n2354, n2351, n2348, n2345, n2342, n2339, n2336, n2333, n2330, n2327, n2324, n2321, n2318, n2315, n2312, n2309, n2306, n2303, n2300, n2297, n2294, n2291, n2288, n2285, n2282, n2279, n2276, n2273, n2270, n2267, n2264, n2261, n2258, n2255, n2252, n2249, n2246, n2243, n2240, n2237, n2234, n2231, n2228, n2225, n2222, n2219, n2216, n2213, n2210};
  /* fplog32.vhdl:1249:4  */
  always @*
    case (n3745)
      512'b10000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b1111111101111100000111111111010101011001;
      512'b01000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b1111111011111100011111111010101011101010;
      512'b00100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b1111111011111100011111111010101011101010;
      512'b00010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b1111111001111101000111101110000101000010;
      512'b00001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b1111111001111101000111101110000101000010;
      512'b00000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b1111110111111101111111010101100101001111;
      512'b00000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b1111110111111101111111010101100101001111;
      512'b00000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b1111110101111111000110101101010001011011;
      512'b00000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b1111110101111111000110101101010001011011;
      512'b00000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b1111110100000000011101110001010000010000;
      512'b00000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b1111110100000000011101110001010000010000;
      512'b00000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b1111110010000010000100011101101001110001;
      512'b00000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b1111110010000010000100011101101001110001;
      512'b00000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b1111110000000011111010101110100111100000;
      512'b00000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b1111110000000011111010101110100111100000;
      512'b00000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b1111101110000110000000100000010100011000;
      512'b00000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b1111101110000110000000100000010100011000;
      512'b00000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b1111101100001000010101101110111100101110;
      512'b00000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b1111101100001000010101101110111100101110;
      512'b00000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b1111101010001010111010010110101110010010;
      512'b00000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b1111101010001010111010010110101110010010;
      512'b00000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b1111101000001101101110010011111000001011;
      512'b00000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b1111101000001101101110010011111000001011;
      512'b00000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b1111100110010000110001100010101010111001;
      512'b00000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b1111100110010000110001100010101010111001;
      512'b00000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b1111100100010100000011111111011000010100;
      512'b00000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b1111100100010100000011111111011000010100;
      512'b00000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b1111100010010111100101100110010011101011;
      512'b00000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b1111100010010111100101100110010011101011;
      512'b00000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b1111100000011011010110010011110001100010;
      512'b00000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b1111100000011011010110010011110001100010;
      512'b00000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b1111011110011111010110000100000111110011;
      512'b00000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b1111011100100011100100110011101101101110;
      512'b00000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b1111011100100011100100110011101101101110;
      512'b00000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b1111011010101000000010011110111011110110;
      512'b00000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b1111011010101000000010011110111011110110;
      512'b00000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b1111011000101100101111000010001100000001;
      512'b00000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b1111011000101100101111000010001100000001;
      512'b00000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b1111010110110001101010011001111001011001;
      512'b00000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b1111010110110001101010011001111001011001;
      512'b00000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b1111010100110110110100100010100000011100;
      512'b00000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b1111010100110110110100100010100000011100;
      512'b00000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b1111010010111100001101011000011110110110;
      512'b00000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b1111010010111100001101011000011110110110;
      512'b00000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b1111010001000001110100111000010011100111;
      512'b00000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b1111001111000111101010111110011110111110;
      512'b00000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b1111001111000111101010111110011110111110;
      512'b00000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b1111001101001101101111100111100010011100;
      512'b00000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b1111001101001101101111100111100010011100;
      512'b00000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b1111001011010100000010110000000000101110;
      512'b00000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b1111001011010100000010110000000000101110;
      512'b00000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b1111001001011010100100010100011101110011;
      512'b00000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b1111001001011010100100010100011101110011;
      512'b00000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b1111000111100001010100010001011110110111;
      512'b00000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b1111000101101000010010100011101010010010;
      512'b00000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b1111000101101000010010100011101010010010;
      512'b00000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b1111000011101111011111000111100111101100;
      512'b00000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b1111000011101111011111000111100111101100;
      512'b00000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b1111000001110110111001111001111111110111;
      512'b00000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b1111000001110110111001111001111111110111;
      512'b00000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b1110111111111110100010110111011100110010;
      512'b00000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b1110111111111110100010110111011100110010;
      512'b00000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b1110111110000110011001111100101001100111;
      512'b00000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b1110111100001110011111000110010010101011;
      512'b00000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b1110111100001110011111000110010010101011;
      512'b00000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b1110111010010110110010010001000101011100;
      512'b00000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b1110111010010110110010010001000101011100;
      512'b00000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b1110111000011111010011011001110000100101;
      512'b00000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b1110111000011111010011011001110000100101;
      512'b00000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b1110110110101000000010011101000011110110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b1110110100110000111111010111110000001010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b1110110100110000111111010111110000001010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b1110110010111010001010000110100111100100;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b1110110010111010001010000110100111100100;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b1110110001000011100010100110011101001110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b1110101111001101001000110100000101011010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b1110101111001101001000110100000101011010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b1110101101010110111100101100010101011110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b1110101101010110111100101100010101011110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b1110101011100000111110001100000011111010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b1110101011100000111110001100000011111010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b1110101001101011001101010000001000010000;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b1110100111110101101001110101011011001001;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b1110100111110101101001110101011011001001;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b1110100110000000010011111000110110010001;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b1110100110000000010011111000110110010001;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b1110100100001011001011010111010100011011;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b1110100010010110010000001101110001011001;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b1110100010010110010000001101110001011001;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b1110100000100001100010011001001010000101;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b1110100000100001100010011001001010000101;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b1110011110101101000001110110011100011000;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b1110011100111000101110100010100111001110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b1110011100111000101110100010100111001110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b1110011011000100101000011010101010100111;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b1110011011000100101000011010101010100111;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b1110011001010000101111011011100111100000;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b1110010111011101000011100010011111111010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b1110010111011101000011100010011111111010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b1110010101101001100100101100010110110101;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b1110010011110110010010110110010000010010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b1110010011110110010010110110010000010010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b1110010010000011001101111101010001001111;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b1110010010000011001101111101010001001111;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b1110010000010000010101111110011111101100;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b1110001110011101101010110111000010100100;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b1110001110011101101010110111000010100100;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b1110001100101011001100100100000001110100;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b1110001100101011001100100100000001110100;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b1110001010111000111011000010100110010011;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b1110001001000110110110001111111001111000;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b1110001001000110110110001111111001111000;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b1110000111010100111110001001000111010101;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b1110000101100011010010101011011010011001;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b1110000101100011010010101011011010011001;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b1110000011110001110011110011111111101111;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b1110000010000000100001100000000100111100;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b1110000010000000100001100000000100111100;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b1110000000001111011011101100111000100100;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b1110000000001111011011101100111000100100;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b1101111110011110100010010111101010000010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b1101111100101101110101011101101001101011;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b1101111100101101110101011101101001101011;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b1101111010111101010100111100001000110010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b1101111001001101000000110000011001011111;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b1101111001001101000000110000011001011111;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b1101110111011100111000110111101110110110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b1101110101101100111101001111011100110010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b1101110101101100111101001111011100110010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b1101110011111101001101110100111000000111;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b1101110010001101101010100101010110100001;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b1101110010001101101010100101010110100001;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b1101110000011110010011011110001110100100;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b1101101110101111001000011100110111101011;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b1101101110101111001000011100110111101011;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b1101101101000000001001011110101010000111;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b1101101011010001010110100000111111000000;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b1101101011010001010110100000111111000000;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b1101101001100010101111100001010000010100;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b1101100111110100010100011100111000110111;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b1101100111110100010100011100111000110111;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b1101100110000110000101010001010100010010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b1101100100011000000001111011111111000011;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b1101100100011000000001111011111111000011;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b1101100010101010001010011010010110011101;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b1101100000111100011110101001111000100110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b1101100000111100011110101001111000100110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b1101011111001110111110101000000100011011;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b1101011101100001101010010010011001101001;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b1101011101100001101010010010011001101001;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b1101011011110100100001100110011000110010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b1101011010000111100100100001100011001011;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b1101011010000111100100100001100011001011;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b1101011000011010110011000001011010111100;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b1101010110101110001101000011100010111100;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b1101010101000001110010100101011110111010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b1101010101000001110010100101011110111010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b1101010011010101100011100100110011010000;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b1101010001101001011111111111000101001101;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b1101010001101001011111111111000101001101;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b1101001111111101100111110001111010110001;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b1101001110010001111010111010111010101011;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b1101001110010001111010111010111010101011;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b1101001100100110011001010111101100011011;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b1101001010111011000011000101111000010001;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b1101001001001111111000000011000111001100;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b1101001001001111111000000011000111001100;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b1101000111100100111000001101000010111101;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b1101000101111010000011100001010110000000;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b1101000101111010000011100001010110000000;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b1101000100001111011001111101101011100010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b1101000010100100111011011111101111011110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b1101000000111010101000000101001110011110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b1101000000111010101000000101001110011110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b1100111111010000011111101011110101111001;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b1100111101100110100010010001010011110011;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b1100111101100110100010010001010011110011;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b1100111011111100101111110011010110111110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b1100111010010011001000001111101110111001;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b1100111000101001101011100100001011101111;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b1100111000101001101011100100001011101111;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b1100110111000000011001101110011110011000;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b1100110101010111010010101100011000010111;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b1100110011101110010110011011101011111101;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b1100110011101110010110011011101011111101;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b1100110010000101100100111010001100000100;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b1100110000011100111110000101101100010011;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b1100101110110100100001111100000000111010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b1100101110110100100001111100000000111010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b1100101101001100010000011010111110111000;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b1100101011100100001001100000011011110000;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b1100101001111100001101001010001101110100;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b1100101001111100001101001010001101110100;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b1100101000010100011011010110001011111110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b1100100110101100110100000010001101110100;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b1100100101000101010111001100001011100000;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b1100100101000101010111001100001011100000;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b1100100011011110000100110001111101111100;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b1100100001110110111100110001011110100101;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b1100100000001111111111001000100111100100;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b1100011110101001001011110101010011101000;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b1100011110101001001011110101010011101000;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b1100011101000010100010110101011110001010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b1100011011011100000100000111000011001011;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b1100011001110101101111100111111111010001;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b1100011001110101101111100111111111010001;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b1100011000001111100101010110001111101100;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b1100010110101001100101001111110010010010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b1100010101000011101111010010100101100000;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b1100010011011110000011011100101000011010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b1100010011011110000011011100101000011010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b1100010001111000100001101011111010101000;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b1100010000010011001001111110011100011100;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b1100001110101101111100010010001110101010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b1100001101001000111000100101010010101111;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b1100001101001000111000100101010010101111;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b1100001011100011111110110101101010101011;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b1100001001111111001111000001011001000101;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b1100001000011010101001000110100001000111;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b1100000110110110001101000011000110100010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b1100000110110110001101000011000110100010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b1100000101010001111010110101001101101001;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b1100000011101101110010011010111011010101;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b1100000010001001110011110010010101000100;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b1100000000100101111110111001100000110100;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b1011111111000010010011101110100101001010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b1011111111000010010011101110100101001010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b1011111101011110110010001111101001010000;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b1011111011111011011010011010110100101100;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b1011111010011000001100001110001111110000;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b1011111000110101000111101000000011001010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b1011111000110101000111101000000011001010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b1011110111010010001100100110011000001110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b1011110101101111011011000111011000110010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b1011110100001100110011001001001111001100;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b1011110010101010010100101010000110010101;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b1011110001000111111111101000001001101010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b1011101111100101110100000001100101000111;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b1011101111100101110100000001100101000111;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b1011101110000011110001110100100101001010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b1011101100100001111000111111010110110010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b1011101011000000001001100000000111011110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b1011101001011110100011010101000101010010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b1011100111111101000110011100011110101100;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b1011100110011011110010110100100010110000;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b1011100110011011110010110100100010110000;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b1011100100111010101000011011100000111110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b1011100011011001100111001111101001011010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b1011100001111000101111001111001100100100;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b1011100000011000000000011000011011011110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b1011011110110111011010101001100111101000;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b1011011101010110111110000001000011000010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b1011011011110110101010011101000000001100;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b1011011011110110101010011101000000001100;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b1011011010010110011111111011110010000010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b1011011000110110011110011011101100000010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b0110011101001000101011111010100001011000;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b0110011010001001010101110000110011110000;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b0110011010001001010101110000110011110000;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b0110010111001010100011010000110001001110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b0110010111001010100011010000110001001110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b0110010100001100010100001101001010000001;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b0110010100001100010100001101001010000001;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b0110010100001100010100001101001010000001;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b0110010001001110101000011000110101110000;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b0110010001001110101000011000110101110000;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b0110001110010001011111100110110011010010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b0110001110010001011111100110110011010010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b0110001011010100111001101010001000101100;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b0110001011010100111001101010001000101100;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b0110001000011000110110010110000011001010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b0110001000011000110110010110000011001010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b0110000101011101010101011101110110110111;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b0110000101011101010101011101110110110111;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b0110000101011101010101011101110110110111;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b0110000010100010010110110100111110111110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b0110000010100010010110110100111110111110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b0101111111100111111010001110111101100000;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b0101111111100111111010001110111101100000;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b0101111100101101111111011111011011010010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b0101111100101101111111011111011011010010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b0101111001110100100110011010000111110100;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b0101111001110100100110011010000111110100;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b0101110110111011101110110010111001010010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b0101110110111011101110110010111001010010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b0101110100000011011000011101101100011010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b0101110100000011011000011101101100011010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b0101110001001011100011001110100100011010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b0101110001001011100011001110100100011010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b0101101110010100001110111001101010111100;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b0101101110010100001110111001101010111100;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b0101101011011101011011010011001111111110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b0101101011011101011011010011001111111110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b0101101000100111001000001111101001110010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b0101101000100111001000001111101001110010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b0101100101110001010101100011010100110100;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b0101100101110001010101100011010100110100;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b0101100010111100000011000010110011101010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b0101100010111100000011000010110011101010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b0101100000000111010000100010101111000010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b0101100000000111010000100010101111000010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b0101011101010010111101110111110101100110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b0101011101010010111101110111110101100110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b0101011010011111001010110110111011111100;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b0101011010011111001010110110111011111100;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b0101010111101011110111010100111100100100;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b0101010111101011110111010100111100100100;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b0101010100111001000011000110110111110000;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b0101010100111001000011000110110111110000;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b0101010010000110101110000001110011100010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b0101010010000110101110000001110011100010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b0101001111010100110111111010111011101010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b0101001111010100110111111010111011101010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b0101001100100011100000100111100001011100;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b0101001100100011100000100111100001011100;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b0101001001110010100111111100111011110011;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b0101001001110010100111111100111011110011;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b0101000111000010001101110000100111000111;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b0101000111000010001101110000100111000111;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b0101000100010010010001111000000101001110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b0101000100010010010001111000000101001110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b0101000001100010110100001000111101011000;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b0101000001100010110100001000111101011000;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b0100111110110011110100011000111100000110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b0100111100000101010010011101110011001101;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b0100111100000101010010011101110011001101;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b0100111001010111001110001101011001101111;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b0100111001010111001110001101011001101111;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b0100110110101001100111011101101011111000;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b0100110110101001100111011101101011111000;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b0100110011111100011110000100101010111011;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b0100110011111100011110000100101010111011;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b0100110001001111110001111000011101001110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b0100110001001111110001111000011101001110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b0100101110100011100010101111001110000100;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b0100101011110111110000011111001101110010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b0100101011110111110000011111001101110010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b0100101001001100011010111110110001100010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b0100101001001100011010111110110001100010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b0100100110100001100010000100010011010100;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b0100100110100001100010000100010011010100;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b0100100011110111000101100110010001111011;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b0100100011110111000101100110010001111011;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b0100100001001101000101011011010000111011;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b0100011110100011100001011001111000100010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b0100011110100011100001011001111000100010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b0100011011111010011001011000110101101010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b0100011011111010011001011000110101101010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b0100011001010001101101001110111001101111;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b0100011001010001101101001110111001101111;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b0100010110101001011100110010111010110100;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b0100010100000001100111111011110011011010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b0100010100000001100111111011110011011010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b0100010001011010001110100000100010100000;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b0100010001011010001110100000100010100000;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b0100001110110011010000011000001011011110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b0100001100001100101101011001110110000110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b0100001100001100101101011001110110000110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b0100001001100110100101011100101110011011;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b0100001001100110100101011100101110011011;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b0100000111000000111000011000000100110110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b0100000111000000111000011000000100110110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b0100000100011011100110000011001101111010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b0100000001110110101110010101100010011011;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b0100000001110110101110010101100010011011;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b0011111111010010010001000110011111010100;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b0011111100101110001110001101100101101000;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b0011111100101110001110001101100101101000;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b0011111010001010100101100010011010011100;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b0011111010001010100101100010011010011100;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b0011110111100111010110111100100110111010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b0011110101000100100010010011111000001001;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b0011110101000100100010010011111000001001;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b0011110010100010000111011111111111001110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b0011110010100010000111011111111111001110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b0011110000000000000110011000110001000111;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b0011101101011110011110110110000110101001;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b0011101101011110011110110110000110101001;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b0011101010111101010000101111111100100000;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b0011101000011100011011111110010011001011;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b0011101000011100011011111110010011001011;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b0011100101111100000000011001001110110110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b0011100101111100000000011001001110110110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b0011100011011011111101111000110111100000;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b0011100000111100010100010101011000110000;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b0011100000111100010100010101011000110000;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b0011011110011101000011100111000001111000;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b0011011011111110001011100110000101110000;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b0011011011111110001011100110000101110000;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b0011011001011111101100001010111010111000;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b0011010111000001100101001101111011001110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b0011010111000001100101001101111011001110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b0011010100100011110110100111100100010110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b0011010010000110100000010000010111001101;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b0011010010000110100000010000010111001101;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b0011001111101001100010000000111000010001;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b0011001101001100111011110001101111010111;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b0011001101001100111011110001101111010111;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b0011001010110000101101011011100111101110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b0011001000010100110110110111001111111010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b0011001000010100110110110111001111111010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b0011000101111001010111111101011001110010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b0011000011011110010000100110111010100010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b0011000011011110010000100110111010100010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b0011000001000011100000101100101010100011;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b0010111110101001001000000111100101011111;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b0010111110101001001000000111100101011111;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b0010111100001111000110110000101010001000;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b0010111001110101011100100000111010100000;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b0010111001110101011100100000111010100000;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b0010110111011100001001010001011011101011;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b0010110101000011001100111011010101111000;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b0010110010101010100111010111110100011000;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b0010110010101010100111010111110100011000;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b0010110000010010011000100000000101100001;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b0010101101111010100000001101011010101000;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b0010101101111010100000001101011010101000;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b0010101011100010111110011001001000000011;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b0010101001001011110010111100100101000100;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b0010100110110100111101110001001011111000;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b0010100110110100111101110001001011111000;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b0010100100011110011110110000011001101000;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b0010100010001000010101110011101110010100;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b0010100010001000010101110011101110010100;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b0010011111110010100010110100101100110010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b0010011101011101000101101100111010110000;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b0010011011000111111110010110000000101011;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b0010011011000111111110010110000000101011;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b0010011000110011001100101001101001110100;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b0010010110011110110000100001100100001101;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b0010010100001010101001110111100000100011;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b0010010100001010101001110111100000100011;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b0010010001110110111000100101010010010100;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b0010001111100011011100100100101111100101;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b0010001101010000010101101111110001001000;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b0010001101010000010101101111110001001000;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b0010001010111101100100000000010010010110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b0010001000101011000111010000010001010000;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b0010000110011000111111011001101110011010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b0010000110011000111111011001101110011010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b0010000100000111001100010110101100111100;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b0010000001110101101110000001010010100100;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b0001111111100100100100010011100111011100;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b0001111111100100100100010011100111011100;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b0001111101010011101111000111110110010000;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b0001111011000011001110011000001100001010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b0001111000110011000001111110111000110000;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b0001110110100011001001110110001110000100;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b0001110110100011001001110110001110000100;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b0001110100010011100101111000100000100010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b0001110010000100010110000000000110111100;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000: n3746 = 40'b0001101111110101011010000111011010100000;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000: n3746 = 40'b0001101101100110110010001000110110101101;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000: n3746 = 40'b0001101101100110110010001000110110101101;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000: n3746 = 40'b0001101011011000011101111110111001011011;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000: n3746 = 40'b0001101001001010011101100100000010110010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000: n3746 = 40'b0001100110111100110000110010110101001101;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000: n3746 = 40'b0001100100101111010111100101110101011001;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000: n3746 = 40'b0001100100101111010111100101110101011001;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000: n3746 = 40'b0001100010100010010001110111101010010010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000: n3746 = 40'b0001100000010101011111100010111101000001;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000: n3746 = 40'b0001011110001001000000100010011000111110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000: n3746 = 40'b0001011011111100110100110000101011101011;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000: n3746 = 40'b0001011001110000111100001000100100110110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000: n3746 = 40'b0001011001110000111100001000100100110110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000: n3746 = 40'b0001010111100101010110100100110110011000;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000: n3746 = 40'b0001010101011010000100000000010100001110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000: n3746 = 40'b0001010011001111000100010101110100100000;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000: n3746 = 40'b0001010001000100010111100000001111011100;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000: n3746 = 40'b0001001110111001111101011010011111010010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000: n3746 = 40'b0001001100101111110101111111100000011000;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000: n3746 = 40'b0001001100101111110101111111100000011000;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000: n3746 = 40'b0001001010100110000001001010010001000111;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000: n3746 = 40'b0001001000011100011110110101110001111000;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000: n3746 = 40'b0001000110010011001110111101000101000110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000: n3746 = 40'b0001000100001010010001011011001111001011;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000: n3746 = 40'b0001000010000001100110001011010110011110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000: n3746 = 40'b0000111111111001001101001000100011010110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000: n3746 = 40'b0000111111111001001101001000100011010110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000: n3746 = 40'b0000111101110001000110001110000000000011;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000: n3746 = 40'b0000111011101001010001010110111000110100;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000: n3746 = 40'b0000111001100001101110011110011011101111;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000: n3746 = 40'b0000110111011010011101011111111000110100;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000: n3746 = 40'b0000110101010011011110010110100001111110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000: n3746 = 40'b0000110011001100110000111101101010111010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000: n3746 = 40'b0000110001000110010101010000101001010000;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000: n3746 = 40'b0000101111000000001011001010110100011011;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000: n3746 = 40'b0000101100111010010010100111100101101010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000: n3746 = 40'b0000101100111010010010100111100101101010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000: n3746 = 40'b0000101010110100101011100010011000000010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000: n3746 = 40'b0000101000101111010101110110101000010111;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000: n3746 = 40'b0000100110101010010001011111110101010001;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000: n3746 = 40'b0000100100100101011110011001011111000111;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000: n3746 = 40'b0000100010100000111100011111001000000000;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000: n3746 = 40'b0000100000011100101011101100010011110100;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000: n3746 = 40'b0000011110011000101011111100101000000101;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000: n3746 = 40'b0000011100010100111101001011101100000101;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000: n3746 = 40'b0000011010010001011111010101001000110001;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000: n3746 = 40'b0000011000001110010010010100101000110010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000: n3746 = 40'b0000010110001011010110000101111000011010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000: n3746 = 40'b0000010100001000101010100100100101100110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000: n3746 = 40'b0000010010000110001111101100011111111011;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000: n3746 = 40'b0000010000000100000101011001011000100101;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000: n3746 = 40'b0000001110000010001011100111000010011001;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000: n3746 = 40'b0000001100000000100010010001010001110001;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000: n3746 = 40'b0000001001111111001001010011111100101101;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000: n3746 = 40'b0000000111111110000000101010111010110001;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000: n3746 = 40'b0000000101111101001000010010000101000110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000: n3746 = 40'b0000000011111100100000000101010110010110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100: n3746 = 40'b0000000001111100001000000000101010101111;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010: n3746 = 40'b1111111111111100000000000000000000000000;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001: n3746 = 40'b1111111111111100000000000000000000000000;
      default: n3746 = 40'bX;
    endcase
  /* fplog32.vhdl:1244:10  */
  always @(posedge clk)
    n3747 <= y0;
  /* fplog32.vhdl:1244:10  */
  always @(posedge clk)
    n3748 <= x;
endmodule

module intadder_27_freq500_uid18
  (input  clk,
   input  [26:0] x,
   input  [26:0] y,
   input  cin,
   output [26:0] r);
  wire cin_0;
  wire cin_0_d1;
  wire cin_0_d2;
  wire cin_0_d3;
  wire cin_0_d4;
  wire cin_0_d5;
  wire cin_0_d6;
  wire [10:0] x_0;
  wire [10:0] x_0_d1;
  wire [10:0] x_0_d2;
  wire [10:0] x_0_d3;
  wire [10:0] y_0;
  wire [10:0] y_0_d1;
  wire [10:0] s_0;
  wire [9:0] r_0;
  wire cin_1;
  wire [17:0] x_1;
  wire [17:0] x_1_d1;
  wire [17:0] x_1_d2;
  wire [17:0] x_1_d3;
  wire [17:0] y_1;
  wire [17:0] y_1_d1;
  wire [17:0] s_1;
  wire [16:0] r_1;
  wire [9:0] n2165;
  wire [10:0] n2167;
  wire [9:0] n2168;
  wire [10:0] n2170;
  wire [10:0] n2171;
  wire [10:0] n2172;
  wire [10:0] n2173;
  wire [9:0] n2174;
  wire n2175;
  wire [16:0] n2176;
  wire [17:0] n2178;
  wire [16:0] n2179;
  wire [17:0] n2181;
  wire [17:0] n2182;
  wire [17:0] n2183;
  wire [17:0] n2184;
  wire [16:0] n2185;
  wire [26:0] n2186;
  reg n2187;
  reg n2188;
  reg n2189;
  reg n2190;
  reg n2191;
  reg n2192;
  reg [10:0] n2193;
  reg [10:0] n2194;
  reg [10:0] n2195;
  reg [10:0] n2196;
  reg [17:0] n2197;
  reg [17:0] n2198;
  reg [17:0] n2199;
  reg [17:0] n2200;
  assign r = n2186; //(module output)
  /* fplog32.vhdl:1152:15  */
  assign cin_0_d1 = n2187; // (signal)
  /* fplog32.vhdl:1152:25  */
  assign cin_0_d2 = n2188; // (signal)
  /* fplog32.vhdl:1152:35  */
  assign cin_0_d3 = n2189; // (signal)
  /* fplog32.vhdl:1152:45  */
  assign cin_0_d4 = n2190; // (signal)
  /* fplog32.vhdl:1152:55  */
  assign cin_0_d5 = n2191; // (signal)
  /* fplog32.vhdl:1152:65  */
  assign cin_0_d6 = n2192; // (signal)
  /* fplog32.vhdl:1154:8  */
  assign x_0 = n2167; // (signal)
  /* fplog32.vhdl:1154:13  */
  assign x_0_d1 = n2193; // (signal)
  /* fplog32.vhdl:1154:21  */
  assign x_0_d2 = n2194; // (signal)
  /* fplog32.vhdl:1154:29  */
  assign x_0_d3 = n2195; // (signal)
  /* fplog32.vhdl:1156:8  */
  assign y_0 = n2170; // (signal)
  /* fplog32.vhdl:1156:13  */
  assign y_0_d1 = n2196; // (signal)
  /* fplog32.vhdl:1158:8  */
  assign s_0 = n2173; // (signal)
  /* fplog32.vhdl:1160:8  */
  assign r_0 = n2174; // (signal)
  /* fplog32.vhdl:1162:8  */
  assign cin_1 = n2175; // (signal)
  /* fplog32.vhdl:1164:8  */
  assign x_1 = n2178; // (signal)
  /* fplog32.vhdl:1164:13  */
  assign x_1_d1 = n2197; // (signal)
  /* fplog32.vhdl:1164:21  */
  assign x_1_d2 = n2198; // (signal)
  /* fplog32.vhdl:1164:29  */
  assign x_1_d3 = n2199; // (signal)
  /* fplog32.vhdl:1166:8  */
  assign y_1 = n2181; // (signal)
  /* fplog32.vhdl:1166:13  */
  assign y_1_d1 = n2200; // (signal)
  /* fplog32.vhdl:1168:8  */
  assign s_1 = n2184; // (signal)
  /* fplog32.vhdl:1170:8  */
  assign r_1 = n2185; // (signal)
  /* fplog32.vhdl:1193:18  */
  assign n2165 = x[9:0]; // extract
  /* fplog32.vhdl:1193:15  */
  assign n2167 = {1'b0, n2165};
  /* fplog32.vhdl:1194:18  */
  assign n2168 = y[9:0]; // extract
  /* fplog32.vhdl:1194:15  */
  assign n2170 = {1'b0, n2168};
  /* fplog32.vhdl:1195:18  */
  assign n2171 = x_0_d3 + y_0_d1;
  /* fplog32.vhdl:1195:27  */
  assign n2172 = {10'b0, cin_0_d6};  //  uext
  /* fplog32.vhdl:1195:27  */
  assign n2173 = n2171 + n2172;
  /* fplog32.vhdl:1196:14  */
  assign n2174 = s_0[9:0]; // extract
  /* fplog32.vhdl:1197:16  */
  assign n2175 = s_0[10]; // extract
  /* fplog32.vhdl:1198:18  */
  assign n2176 = x[26:10]; // extract
  /* fplog32.vhdl:1198:15  */
  assign n2178 = {1'b0, n2176};
  /* fplog32.vhdl:1199:18  */
  assign n2179 = y[26:10]; // extract
  /* fplog32.vhdl:1199:15  */
  assign n2181 = {1'b0, n2179};
  /* fplog32.vhdl:1200:18  */
  assign n2182 = x_1_d3 + y_1_d1;
  /* fplog32.vhdl:1200:27  */
  assign n2183 = {17'b0, cin_1};  //  uext
  /* fplog32.vhdl:1200:27  */
  assign n2184 = n2182 + n2183;
  /* fplog32.vhdl:1201:14  */
  assign n2185 = s_1[16:0]; // extract
  /* fplog32.vhdl:1202:13  */
  assign n2186 = {r_1, r_0};
  /* fplog32.vhdl:1175:10  */
  always @(posedge clk)
    n2187 <= cin_0;
  /* fplog32.vhdl:1175:10  */
  always @(posedge clk)
    n2188 <= cin_0_d1;
  /* fplog32.vhdl:1175:10  */
  always @(posedge clk)
    n2189 <= cin_0_d2;
  /* fplog32.vhdl:1175:10  */
  always @(posedge clk)
    n2190 <= cin_0_d3;
  /* fplog32.vhdl:1175:10  */
  always @(posedge clk)
    n2191 <= cin_0_d4;
  /* fplog32.vhdl:1175:10  */
  always @(posedge clk)
    n2192 <= cin_0_d5;
  /* fplog32.vhdl:1175:10  */
  always @(posedge clk)
    n2193 <= x_0;
  /* fplog32.vhdl:1175:10  */
  always @(posedge clk)
    n2194 <= x_0_d1;
  /* fplog32.vhdl:1175:10  */
  always @(posedge clk)
    n2195 <= x_0_d2;
  /* fplog32.vhdl:1175:10  */
  always @(posedge clk)
    n2196 <= y_0;
  /* fplog32.vhdl:1175:10  */
  always @(posedge clk)
    n2197 <= x_1;
  /* fplog32.vhdl:1175:10  */
  always @(posedge clk)
    n2198 <= x_1_d1;
  /* fplog32.vhdl:1175:10  */
  always @(posedge clk)
    n2199 <= x_1_d2;
  /* fplog32.vhdl:1175:10  */
  always @(posedge clk)
    n2200 <= y_1;
endmodule

module intadder_27_freq500_uid15
  (input  clk,
   input  [26:0] x,
   input  [26:0] y,
   input  cin,
   output [26:0] r);
  wire cin_1;
  wire cin_1_d1;
  wire cin_1_d2;
  wire cin_1_d3;
  wire [27:0] x_1;
  wire [27:0] x_1_d1;
  wire [27:0] y_1;
  wire [27:0] y_1_d1;
  wire [27:0] s_1;
  wire [26:0] r_1;
  wire [27:0] n2134;
  wire [27:0] n2136;
  wire [27:0] n2137;
  wire [27:0] n2138;
  wire [27:0] n2139;
  wire [26:0] n2140;
  reg n2141;
  reg n2142;
  reg n2143;
  reg [27:0] n2144;
  reg [27:0] n2145;
  assign r = r_1; //(module output)
  /* fplog32.vhdl:1091:15  */
  assign cin_1_d1 = n2141; // (signal)
  /* fplog32.vhdl:1091:25  */
  assign cin_1_d2 = n2142; // (signal)
  /* fplog32.vhdl:1091:35  */
  assign cin_1_d3 = n2143; // (signal)
  /* fplog32.vhdl:1093:8  */
  assign x_1 = n2134; // (signal)
  /* fplog32.vhdl:1093:13  */
  assign x_1_d1 = n2144; // (signal)
  /* fplog32.vhdl:1095:8  */
  assign y_1 = n2136; // (signal)
  /* fplog32.vhdl:1095:13  */
  assign y_1_d1 = n2145; // (signal)
  /* fplog32.vhdl:1097:8  */
  assign s_1 = n2139; // (signal)
  /* fplog32.vhdl:1099:8  */
  assign r_1 = n2140; // (signal)
  /* fplog32.vhdl:1113:15  */
  assign n2134 = {1'b0, x};
  /* fplog32.vhdl:1114:15  */
  assign n2136 = {1'b0, y};
  /* fplog32.vhdl:1115:18  */
  assign n2137 = x_1_d1 + y_1_d1;
  /* fplog32.vhdl:1115:27  */
  assign n2138 = {27'b0, cin_1_d3};  //  uext
  /* fplog32.vhdl:1115:27  */
  assign n2139 = n2137 + n2138;
  /* fplog32.vhdl:1116:14  */
  assign n2140 = s_1[26:0]; // extract
  /* fplog32.vhdl:1104:10  */
  always @(posedge clk)
    n2141 <= cin_1;
  /* fplog32.vhdl:1104:10  */
  always @(posedge clk)
    n2142 <= cin_1_d1;
  /* fplog32.vhdl:1104:10  */
  always @(posedge clk)
    n2143 <= cin_1_d2;
  /* fplog32.vhdl:1104:10  */
  always @(posedge clk)
    n2144 <= x_1;
  /* fplog32.vhdl:1104:10  */
  always @(posedge clk)
    n2145 <= y_1;
endmodule

module intadder_27_freq500_uid12
  (input  clk,
   input  [26:0] x,
   input  [26:0] y,
   input  cin,
   output [26:0] r);
  wire cin_1;
  wire cin_1_d1;
  wire cin_1_d2;
  wire [27:0] x_1;
  wire [27:0] x_1_d1;
  wire [27:0] y_1;
  wire [27:0] y_1_d1;
  wire [27:0] s_1;
  wire [26:0] r_1;
  wire [27:0] n2112;
  wire [27:0] n2114;
  wire [27:0] n2115;
  wire [27:0] n2116;
  wire [27:0] n2117;
  wire [26:0] n2118;
  reg n2119;
  reg n2120;
  reg [27:0] n2121;
  reg [27:0] n2122;
  assign r = r_1; //(module output)
  /* fplog32.vhdl:1031:15  */
  assign cin_1_d1 = n2119; // (signal)
  /* fplog32.vhdl:1031:25  */
  assign cin_1_d2 = n2120; // (signal)
  /* fplog32.vhdl:1033:8  */
  assign x_1 = n2112; // (signal)
  /* fplog32.vhdl:1033:13  */
  assign x_1_d1 = n2121; // (signal)
  /* fplog32.vhdl:1035:8  */
  assign y_1 = n2114; // (signal)
  /* fplog32.vhdl:1035:13  */
  assign y_1_d1 = n2122; // (signal)
  /* fplog32.vhdl:1037:8  */
  assign s_1 = n2117; // (signal)
  /* fplog32.vhdl:1039:8  */
  assign r_1 = n2118; // (signal)
  /* fplog32.vhdl:1052:15  */
  assign n2112 = {1'b0, x};
  /* fplog32.vhdl:1053:15  */
  assign n2114 = {1'b0, y};
  /* fplog32.vhdl:1054:18  */
  assign n2115 = x_1_d1 + y_1_d1;
  /* fplog32.vhdl:1054:27  */
  assign n2116 = {27'b0, cin_1_d2};  //  uext
  /* fplog32.vhdl:1054:27  */
  assign n2117 = n2115 + n2116;
  /* fplog32.vhdl:1055:14  */
  assign n2118 = s_1[26:0]; // extract
  /* fplog32.vhdl:1044:10  */
  always @(posedge clk)
    n2119 <= cin_1;
  /* fplog32.vhdl:1044:10  */
  always @(posedge clk)
    n2120 <= cin_1_d1;
  /* fplog32.vhdl:1044:10  */
  always @(posedge clk)
    n2121 <= x_1;
  /* fplog32.vhdl:1044:10  */
  always @(posedge clk)
    n2122 <= y_1;
endmodule

module inva0table_freq500_uid8
  (input  [8:0] x,
   output [9:0] y);
  wire [9:0] y0;
  wire [9:0] y1;
  wire n565;
  wire n568;
  wire n571;
  wire n574;
  wire n577;
  wire n580;
  wire n583;
  wire n586;
  wire n589;
  wire n592;
  wire n595;
  wire n598;
  wire n601;
  wire n604;
  wire n607;
  wire n610;
  wire n613;
  wire n616;
  wire n619;
  wire n622;
  wire n625;
  wire n628;
  wire n631;
  wire n634;
  wire n637;
  wire n640;
  wire n643;
  wire n646;
  wire n649;
  wire n652;
  wire n655;
  wire n658;
  wire n661;
  wire n664;
  wire n667;
  wire n670;
  wire n673;
  wire n676;
  wire n679;
  wire n682;
  wire n685;
  wire n688;
  wire n691;
  wire n694;
  wire n697;
  wire n700;
  wire n703;
  wire n706;
  wire n709;
  wire n712;
  wire n715;
  wire n718;
  wire n721;
  wire n724;
  wire n727;
  wire n730;
  wire n733;
  wire n736;
  wire n739;
  wire n742;
  wire n745;
  wire n748;
  wire n751;
  wire n754;
  wire n757;
  wire n760;
  wire n763;
  wire n766;
  wire n769;
  wire n772;
  wire n775;
  wire n778;
  wire n781;
  wire n784;
  wire n787;
  wire n790;
  wire n793;
  wire n796;
  wire n799;
  wire n802;
  wire n805;
  wire n808;
  wire n811;
  wire n814;
  wire n817;
  wire n820;
  wire n823;
  wire n826;
  wire n829;
  wire n832;
  wire n835;
  wire n838;
  wire n841;
  wire n844;
  wire n847;
  wire n850;
  wire n853;
  wire n856;
  wire n859;
  wire n862;
  wire n865;
  wire n868;
  wire n871;
  wire n874;
  wire n877;
  wire n880;
  wire n883;
  wire n886;
  wire n889;
  wire n892;
  wire n895;
  wire n898;
  wire n901;
  wire n904;
  wire n907;
  wire n910;
  wire n913;
  wire n916;
  wire n919;
  wire n922;
  wire n925;
  wire n928;
  wire n931;
  wire n934;
  wire n937;
  wire n940;
  wire n943;
  wire n946;
  wire n949;
  wire n952;
  wire n955;
  wire n958;
  wire n961;
  wire n964;
  wire n967;
  wire n970;
  wire n973;
  wire n976;
  wire n979;
  wire n982;
  wire n985;
  wire n988;
  wire n991;
  wire n994;
  wire n997;
  wire n1000;
  wire n1003;
  wire n1006;
  wire n1009;
  wire n1012;
  wire n1015;
  wire n1018;
  wire n1021;
  wire n1024;
  wire n1027;
  wire n1030;
  wire n1033;
  wire n1036;
  wire n1039;
  wire n1042;
  wire n1045;
  wire n1048;
  wire n1051;
  wire n1054;
  wire n1057;
  wire n1060;
  wire n1063;
  wire n1066;
  wire n1069;
  wire n1072;
  wire n1075;
  wire n1078;
  wire n1081;
  wire n1084;
  wire n1087;
  wire n1090;
  wire n1093;
  wire n1096;
  wire n1099;
  wire n1102;
  wire n1105;
  wire n1108;
  wire n1111;
  wire n1114;
  wire n1117;
  wire n1120;
  wire n1123;
  wire n1126;
  wire n1129;
  wire n1132;
  wire n1135;
  wire n1138;
  wire n1141;
  wire n1144;
  wire n1147;
  wire n1150;
  wire n1153;
  wire n1156;
  wire n1159;
  wire n1162;
  wire n1165;
  wire n1168;
  wire n1171;
  wire n1174;
  wire n1177;
  wire n1180;
  wire n1183;
  wire n1186;
  wire n1189;
  wire n1192;
  wire n1195;
  wire n1198;
  wire n1201;
  wire n1204;
  wire n1207;
  wire n1210;
  wire n1213;
  wire n1216;
  wire n1219;
  wire n1222;
  wire n1225;
  wire n1228;
  wire n1231;
  wire n1234;
  wire n1237;
  wire n1240;
  wire n1243;
  wire n1246;
  wire n1249;
  wire n1252;
  wire n1255;
  wire n1258;
  wire n1261;
  wire n1264;
  wire n1267;
  wire n1270;
  wire n1273;
  wire n1276;
  wire n1279;
  wire n1282;
  wire n1285;
  wire n1288;
  wire n1291;
  wire n1294;
  wire n1297;
  wire n1300;
  wire n1303;
  wire n1306;
  wire n1309;
  wire n1312;
  wire n1315;
  wire n1318;
  wire n1321;
  wire n1324;
  wire n1327;
  wire n1330;
  wire n1333;
  wire n1336;
  wire n1339;
  wire n1342;
  wire n1345;
  wire n1348;
  wire n1351;
  wire n1354;
  wire n1357;
  wire n1360;
  wire n1363;
  wire n1366;
  wire n1369;
  wire n1372;
  wire n1375;
  wire n1378;
  wire n1381;
  wire n1384;
  wire n1387;
  wire n1390;
  wire n1393;
  wire n1396;
  wire n1399;
  wire n1402;
  wire n1405;
  wire n1408;
  wire n1411;
  wire n1414;
  wire n1417;
  wire n1420;
  wire n1423;
  wire n1426;
  wire n1429;
  wire n1432;
  wire n1435;
  wire n1438;
  wire n1441;
  wire n1444;
  wire n1447;
  wire n1450;
  wire n1453;
  wire n1456;
  wire n1459;
  wire n1462;
  wire n1465;
  wire n1468;
  wire n1471;
  wire n1474;
  wire n1477;
  wire n1480;
  wire n1483;
  wire n1486;
  wire n1489;
  wire n1492;
  wire n1495;
  wire n1498;
  wire n1501;
  wire n1504;
  wire n1507;
  wire n1510;
  wire n1513;
  wire n1516;
  wire n1519;
  wire n1522;
  wire n1525;
  wire n1528;
  wire n1531;
  wire n1534;
  wire n1537;
  wire n1540;
  wire n1543;
  wire n1546;
  wire n1549;
  wire n1552;
  wire n1555;
  wire n1558;
  wire n1561;
  wire n1564;
  wire n1567;
  wire n1570;
  wire n1573;
  wire n1576;
  wire n1579;
  wire n1582;
  wire n1585;
  wire n1588;
  wire n1591;
  wire n1594;
  wire n1597;
  wire n1600;
  wire n1603;
  wire n1606;
  wire n1609;
  wire n1612;
  wire n1615;
  wire n1618;
  wire n1621;
  wire n1624;
  wire n1627;
  wire n1630;
  wire n1633;
  wire n1636;
  wire n1639;
  wire n1642;
  wire n1645;
  wire n1648;
  wire n1651;
  wire n1654;
  wire n1657;
  wire n1660;
  wire n1663;
  wire n1666;
  wire n1669;
  wire n1672;
  wire n1675;
  wire n1678;
  wire n1681;
  wire n1684;
  wire n1687;
  wire n1690;
  wire n1693;
  wire n1696;
  wire n1699;
  wire n1702;
  wire n1705;
  wire n1708;
  wire n1711;
  wire n1714;
  wire n1717;
  wire n1720;
  wire n1723;
  wire n1726;
  wire n1729;
  wire n1732;
  wire n1735;
  wire n1738;
  wire n1741;
  wire n1744;
  wire n1747;
  wire n1750;
  wire n1753;
  wire n1756;
  wire n1759;
  wire n1762;
  wire n1765;
  wire n1768;
  wire n1771;
  wire n1774;
  wire n1777;
  wire n1780;
  wire n1783;
  wire n1786;
  wire n1789;
  wire n1792;
  wire n1795;
  wire n1798;
  wire n1801;
  wire n1804;
  wire n1807;
  wire n1810;
  wire n1813;
  wire n1816;
  wire n1819;
  wire n1822;
  wire n1825;
  wire n1828;
  wire n1831;
  wire n1834;
  wire n1837;
  wire n1840;
  wire n1843;
  wire n1846;
  wire n1849;
  wire n1852;
  wire n1855;
  wire n1858;
  wire n1861;
  wire n1864;
  wire n1867;
  wire n1870;
  wire n1873;
  wire n1876;
  wire n1879;
  wire n1882;
  wire n1885;
  wire n1888;
  wire n1891;
  wire n1894;
  wire n1897;
  wire n1900;
  wire n1903;
  wire n1906;
  wire n1909;
  wire n1912;
  wire n1915;
  wire n1918;
  wire n1921;
  wire n1924;
  wire n1927;
  wire n1930;
  wire n1933;
  wire n1936;
  wire n1939;
  wire n1942;
  wire n1945;
  wire n1948;
  wire n1951;
  wire n1954;
  wire n1957;
  wire n1960;
  wire n1963;
  wire n1966;
  wire n1969;
  wire n1972;
  wire n1975;
  wire n1978;
  wire n1981;
  wire n1984;
  wire n1987;
  wire n1990;
  wire n1993;
  wire n1996;
  wire n1999;
  wire n2002;
  wire n2005;
  wire n2008;
  wire n2011;
  wire n2014;
  wire n2017;
  wire n2020;
  wire n2023;
  wire n2026;
  wire n2029;
  wire n2032;
  wire n2035;
  wire n2038;
  wire n2041;
  wire n2044;
  wire n2047;
  wire n2050;
  wire n2053;
  wire n2056;
  wire n2059;
  wire n2062;
  wire n2065;
  wire n2068;
  wire n2071;
  wire n2074;
  wire n2077;
  wire n2080;
  wire n2083;
  wire n2086;
  wire n2089;
  wire n2092;
  wire n2095;
  wire n2098;
  wire [511:0] n2100;
  reg [9:0] n2101;
  assign y = y1; //(module output)
  /* fplog32.vhdl:30:8  */
  assign y0 = n2101; // (signal)
  /* fplog32.vhdl:32:8  */
  assign y1 = y0; // (signal)
  /* fplog32.vhdl:36:20  */
  assign n565 = x == 9'b000000000;
  /* fplog32.vhdl:37:20  */
  assign n568 = x == 9'b000000001;
  /* fplog32.vhdl:38:20  */
  assign n571 = x == 9'b000000010;
  /* fplog32.vhdl:39:20  */
  assign n574 = x == 9'b000000011;
  /* fplog32.vhdl:40:20  */
  assign n577 = x == 9'b000000100;
  /* fplog32.vhdl:41:20  */
  assign n580 = x == 9'b000000101;
  /* fplog32.vhdl:42:20  */
  assign n583 = x == 9'b000000110;
  /* fplog32.vhdl:43:20  */
  assign n586 = x == 9'b000000111;
  /* fplog32.vhdl:44:20  */
  assign n589 = x == 9'b000001000;
  /* fplog32.vhdl:45:20  */
  assign n592 = x == 9'b000001001;
  /* fplog32.vhdl:46:20  */
  assign n595 = x == 9'b000001010;
  /* fplog32.vhdl:47:20  */
  assign n598 = x == 9'b000001011;
  /* fplog32.vhdl:48:20  */
  assign n601 = x == 9'b000001100;
  /* fplog32.vhdl:49:20  */
  assign n604 = x == 9'b000001101;
  /* fplog32.vhdl:50:20  */
  assign n607 = x == 9'b000001110;
  /* fplog32.vhdl:51:20  */
  assign n610 = x == 9'b000001111;
  /* fplog32.vhdl:52:20  */
  assign n613 = x == 9'b000010000;
  /* fplog32.vhdl:53:20  */
  assign n616 = x == 9'b000010001;
  /* fplog32.vhdl:54:20  */
  assign n619 = x == 9'b000010010;
  /* fplog32.vhdl:55:20  */
  assign n622 = x == 9'b000010011;
  /* fplog32.vhdl:56:20  */
  assign n625 = x == 9'b000010100;
  /* fplog32.vhdl:57:20  */
  assign n628 = x == 9'b000010101;
  /* fplog32.vhdl:58:20  */
  assign n631 = x == 9'b000010110;
  /* fplog32.vhdl:59:20  */
  assign n634 = x == 9'b000010111;
  /* fplog32.vhdl:60:20  */
  assign n637 = x == 9'b000011000;
  /* fplog32.vhdl:61:20  */
  assign n640 = x == 9'b000011001;
  /* fplog32.vhdl:62:20  */
  assign n643 = x == 9'b000011010;
  /* fplog32.vhdl:63:20  */
  assign n646 = x == 9'b000011011;
  /* fplog32.vhdl:64:20  */
  assign n649 = x == 9'b000011100;
  /* fplog32.vhdl:65:20  */
  assign n652 = x == 9'b000011101;
  /* fplog32.vhdl:66:20  */
  assign n655 = x == 9'b000011110;
  /* fplog32.vhdl:67:20  */
  assign n658 = x == 9'b000011111;
  /* fplog32.vhdl:68:20  */
  assign n661 = x == 9'b000100000;
  /* fplog32.vhdl:69:20  */
  assign n664 = x == 9'b000100001;
  /* fplog32.vhdl:70:20  */
  assign n667 = x == 9'b000100010;
  /* fplog32.vhdl:71:20  */
  assign n670 = x == 9'b000100011;
  /* fplog32.vhdl:72:20  */
  assign n673 = x == 9'b000100100;
  /* fplog32.vhdl:73:20  */
  assign n676 = x == 9'b000100101;
  /* fplog32.vhdl:74:20  */
  assign n679 = x == 9'b000100110;
  /* fplog32.vhdl:75:20  */
  assign n682 = x == 9'b000100111;
  /* fplog32.vhdl:76:20  */
  assign n685 = x == 9'b000101000;
  /* fplog32.vhdl:77:20  */
  assign n688 = x == 9'b000101001;
  /* fplog32.vhdl:78:20  */
  assign n691 = x == 9'b000101010;
  /* fplog32.vhdl:79:20  */
  assign n694 = x == 9'b000101011;
  /* fplog32.vhdl:80:20  */
  assign n697 = x == 9'b000101100;
  /* fplog32.vhdl:81:20  */
  assign n700 = x == 9'b000101101;
  /* fplog32.vhdl:82:20  */
  assign n703 = x == 9'b000101110;
  /* fplog32.vhdl:83:20  */
  assign n706 = x == 9'b000101111;
  /* fplog32.vhdl:84:20  */
  assign n709 = x == 9'b000110000;
  /* fplog32.vhdl:85:20  */
  assign n712 = x == 9'b000110001;
  /* fplog32.vhdl:86:20  */
  assign n715 = x == 9'b000110010;
  /* fplog32.vhdl:87:20  */
  assign n718 = x == 9'b000110011;
  /* fplog32.vhdl:88:20  */
  assign n721 = x == 9'b000110100;
  /* fplog32.vhdl:89:20  */
  assign n724 = x == 9'b000110101;
  /* fplog32.vhdl:90:20  */
  assign n727 = x == 9'b000110110;
  /* fplog32.vhdl:91:20  */
  assign n730 = x == 9'b000110111;
  /* fplog32.vhdl:92:20  */
  assign n733 = x == 9'b000111000;
  /* fplog32.vhdl:93:20  */
  assign n736 = x == 9'b000111001;
  /* fplog32.vhdl:94:20  */
  assign n739 = x == 9'b000111010;
  /* fplog32.vhdl:95:20  */
  assign n742 = x == 9'b000111011;
  /* fplog32.vhdl:96:20  */
  assign n745 = x == 9'b000111100;
  /* fplog32.vhdl:97:20  */
  assign n748 = x == 9'b000111101;
  /* fplog32.vhdl:98:20  */
  assign n751 = x == 9'b000111110;
  /* fplog32.vhdl:99:20  */
  assign n754 = x == 9'b000111111;
  /* fplog32.vhdl:100:20  */
  assign n757 = x == 9'b001000000;
  /* fplog32.vhdl:101:20  */
  assign n760 = x == 9'b001000001;
  /* fplog32.vhdl:102:20  */
  assign n763 = x == 9'b001000010;
  /* fplog32.vhdl:103:20  */
  assign n766 = x == 9'b001000011;
  /* fplog32.vhdl:104:20  */
  assign n769 = x == 9'b001000100;
  /* fplog32.vhdl:105:20  */
  assign n772 = x == 9'b001000101;
  /* fplog32.vhdl:106:20  */
  assign n775 = x == 9'b001000110;
  /* fplog32.vhdl:107:20  */
  assign n778 = x == 9'b001000111;
  /* fplog32.vhdl:108:20  */
  assign n781 = x == 9'b001001000;
  /* fplog32.vhdl:109:20  */
  assign n784 = x == 9'b001001001;
  /* fplog32.vhdl:110:20  */
  assign n787 = x == 9'b001001010;
  /* fplog32.vhdl:111:20  */
  assign n790 = x == 9'b001001011;
  /* fplog32.vhdl:112:20  */
  assign n793 = x == 9'b001001100;
  /* fplog32.vhdl:113:20  */
  assign n796 = x == 9'b001001101;
  /* fplog32.vhdl:114:20  */
  assign n799 = x == 9'b001001110;
  /* fplog32.vhdl:115:20  */
  assign n802 = x == 9'b001001111;
  /* fplog32.vhdl:116:20  */
  assign n805 = x == 9'b001010000;
  /* fplog32.vhdl:117:20  */
  assign n808 = x == 9'b001010001;
  /* fplog32.vhdl:118:20  */
  assign n811 = x == 9'b001010010;
  /* fplog32.vhdl:119:20  */
  assign n814 = x == 9'b001010011;
  /* fplog32.vhdl:120:20  */
  assign n817 = x == 9'b001010100;
  /* fplog32.vhdl:121:20  */
  assign n820 = x == 9'b001010101;
  /* fplog32.vhdl:122:20  */
  assign n823 = x == 9'b001010110;
  /* fplog32.vhdl:123:20  */
  assign n826 = x == 9'b001010111;
  /* fplog32.vhdl:124:20  */
  assign n829 = x == 9'b001011000;
  /* fplog32.vhdl:125:20  */
  assign n832 = x == 9'b001011001;
  /* fplog32.vhdl:126:20  */
  assign n835 = x == 9'b001011010;
  /* fplog32.vhdl:127:20  */
  assign n838 = x == 9'b001011011;
  /* fplog32.vhdl:128:20  */
  assign n841 = x == 9'b001011100;
  /* fplog32.vhdl:129:20  */
  assign n844 = x == 9'b001011101;
  /* fplog32.vhdl:130:20  */
  assign n847 = x == 9'b001011110;
  /* fplog32.vhdl:131:20  */
  assign n850 = x == 9'b001011111;
  /* fplog32.vhdl:132:20  */
  assign n853 = x == 9'b001100000;
  /* fplog32.vhdl:133:20  */
  assign n856 = x == 9'b001100001;
  /* fplog32.vhdl:134:20  */
  assign n859 = x == 9'b001100010;
  /* fplog32.vhdl:135:20  */
  assign n862 = x == 9'b001100011;
  /* fplog32.vhdl:136:20  */
  assign n865 = x == 9'b001100100;
  /* fplog32.vhdl:137:20  */
  assign n868 = x == 9'b001100101;
  /* fplog32.vhdl:138:20  */
  assign n871 = x == 9'b001100110;
  /* fplog32.vhdl:139:20  */
  assign n874 = x == 9'b001100111;
  /* fplog32.vhdl:140:20  */
  assign n877 = x == 9'b001101000;
  /* fplog32.vhdl:141:20  */
  assign n880 = x == 9'b001101001;
  /* fplog32.vhdl:142:20  */
  assign n883 = x == 9'b001101010;
  /* fplog32.vhdl:143:20  */
  assign n886 = x == 9'b001101011;
  /* fplog32.vhdl:144:20  */
  assign n889 = x == 9'b001101100;
  /* fplog32.vhdl:145:20  */
  assign n892 = x == 9'b001101101;
  /* fplog32.vhdl:146:20  */
  assign n895 = x == 9'b001101110;
  /* fplog32.vhdl:147:20  */
  assign n898 = x == 9'b001101111;
  /* fplog32.vhdl:148:20  */
  assign n901 = x == 9'b001110000;
  /* fplog32.vhdl:149:20  */
  assign n904 = x == 9'b001110001;
  /* fplog32.vhdl:150:20  */
  assign n907 = x == 9'b001110010;
  /* fplog32.vhdl:151:20  */
  assign n910 = x == 9'b001110011;
  /* fplog32.vhdl:152:20  */
  assign n913 = x == 9'b001110100;
  /* fplog32.vhdl:153:20  */
  assign n916 = x == 9'b001110101;
  /* fplog32.vhdl:154:20  */
  assign n919 = x == 9'b001110110;
  /* fplog32.vhdl:155:20  */
  assign n922 = x == 9'b001110111;
  /* fplog32.vhdl:156:20  */
  assign n925 = x == 9'b001111000;
  /* fplog32.vhdl:157:20  */
  assign n928 = x == 9'b001111001;
  /* fplog32.vhdl:158:20  */
  assign n931 = x == 9'b001111010;
  /* fplog32.vhdl:159:20  */
  assign n934 = x == 9'b001111011;
  /* fplog32.vhdl:160:20  */
  assign n937 = x == 9'b001111100;
  /* fplog32.vhdl:161:20  */
  assign n940 = x == 9'b001111101;
  /* fplog32.vhdl:162:20  */
  assign n943 = x == 9'b001111110;
  /* fplog32.vhdl:163:20  */
  assign n946 = x == 9'b001111111;
  /* fplog32.vhdl:164:20  */
  assign n949 = x == 9'b010000000;
  /* fplog32.vhdl:165:20  */
  assign n952 = x == 9'b010000001;
  /* fplog32.vhdl:166:20  */
  assign n955 = x == 9'b010000010;
  /* fplog32.vhdl:167:20  */
  assign n958 = x == 9'b010000011;
  /* fplog32.vhdl:168:20  */
  assign n961 = x == 9'b010000100;
  /* fplog32.vhdl:169:20  */
  assign n964 = x == 9'b010000101;
  /* fplog32.vhdl:170:20  */
  assign n967 = x == 9'b010000110;
  /* fplog32.vhdl:171:20  */
  assign n970 = x == 9'b010000111;
  /* fplog32.vhdl:172:20  */
  assign n973 = x == 9'b010001000;
  /* fplog32.vhdl:173:20  */
  assign n976 = x == 9'b010001001;
  /* fplog32.vhdl:174:20  */
  assign n979 = x == 9'b010001010;
  /* fplog32.vhdl:175:20  */
  assign n982 = x == 9'b010001011;
  /* fplog32.vhdl:176:20  */
  assign n985 = x == 9'b010001100;
  /* fplog32.vhdl:177:20  */
  assign n988 = x == 9'b010001101;
  /* fplog32.vhdl:178:20  */
  assign n991 = x == 9'b010001110;
  /* fplog32.vhdl:179:20  */
  assign n994 = x == 9'b010001111;
  /* fplog32.vhdl:180:20  */
  assign n997 = x == 9'b010010000;
  /* fplog32.vhdl:181:20  */
  assign n1000 = x == 9'b010010001;
  /* fplog32.vhdl:182:20  */
  assign n1003 = x == 9'b010010010;
  /* fplog32.vhdl:183:20  */
  assign n1006 = x == 9'b010010011;
  /* fplog32.vhdl:184:20  */
  assign n1009 = x == 9'b010010100;
  /* fplog32.vhdl:185:20  */
  assign n1012 = x == 9'b010010101;
  /* fplog32.vhdl:186:20  */
  assign n1015 = x == 9'b010010110;
  /* fplog32.vhdl:187:20  */
  assign n1018 = x == 9'b010010111;
  /* fplog32.vhdl:188:20  */
  assign n1021 = x == 9'b010011000;
  /* fplog32.vhdl:189:20  */
  assign n1024 = x == 9'b010011001;
  /* fplog32.vhdl:190:20  */
  assign n1027 = x == 9'b010011010;
  /* fplog32.vhdl:191:20  */
  assign n1030 = x == 9'b010011011;
  /* fplog32.vhdl:192:20  */
  assign n1033 = x == 9'b010011100;
  /* fplog32.vhdl:193:20  */
  assign n1036 = x == 9'b010011101;
  /* fplog32.vhdl:194:20  */
  assign n1039 = x == 9'b010011110;
  /* fplog32.vhdl:195:20  */
  assign n1042 = x == 9'b010011111;
  /* fplog32.vhdl:196:20  */
  assign n1045 = x == 9'b010100000;
  /* fplog32.vhdl:197:20  */
  assign n1048 = x == 9'b010100001;
  /* fplog32.vhdl:198:20  */
  assign n1051 = x == 9'b010100010;
  /* fplog32.vhdl:199:20  */
  assign n1054 = x == 9'b010100011;
  /* fplog32.vhdl:200:20  */
  assign n1057 = x == 9'b010100100;
  /* fplog32.vhdl:201:20  */
  assign n1060 = x == 9'b010100101;
  /* fplog32.vhdl:202:20  */
  assign n1063 = x == 9'b010100110;
  /* fplog32.vhdl:203:20  */
  assign n1066 = x == 9'b010100111;
  /* fplog32.vhdl:204:20  */
  assign n1069 = x == 9'b010101000;
  /* fplog32.vhdl:205:20  */
  assign n1072 = x == 9'b010101001;
  /* fplog32.vhdl:206:20  */
  assign n1075 = x == 9'b010101010;
  /* fplog32.vhdl:207:20  */
  assign n1078 = x == 9'b010101011;
  /* fplog32.vhdl:208:20  */
  assign n1081 = x == 9'b010101100;
  /* fplog32.vhdl:209:20  */
  assign n1084 = x == 9'b010101101;
  /* fplog32.vhdl:210:20  */
  assign n1087 = x == 9'b010101110;
  /* fplog32.vhdl:211:20  */
  assign n1090 = x == 9'b010101111;
  /* fplog32.vhdl:212:20  */
  assign n1093 = x == 9'b010110000;
  /* fplog32.vhdl:213:20  */
  assign n1096 = x == 9'b010110001;
  /* fplog32.vhdl:214:20  */
  assign n1099 = x == 9'b010110010;
  /* fplog32.vhdl:215:20  */
  assign n1102 = x == 9'b010110011;
  /* fplog32.vhdl:216:20  */
  assign n1105 = x == 9'b010110100;
  /* fplog32.vhdl:217:20  */
  assign n1108 = x == 9'b010110101;
  /* fplog32.vhdl:218:20  */
  assign n1111 = x == 9'b010110110;
  /* fplog32.vhdl:219:20  */
  assign n1114 = x == 9'b010110111;
  /* fplog32.vhdl:220:20  */
  assign n1117 = x == 9'b010111000;
  /* fplog32.vhdl:221:20  */
  assign n1120 = x == 9'b010111001;
  /* fplog32.vhdl:222:20  */
  assign n1123 = x == 9'b010111010;
  /* fplog32.vhdl:223:20  */
  assign n1126 = x == 9'b010111011;
  /* fplog32.vhdl:224:20  */
  assign n1129 = x == 9'b010111100;
  /* fplog32.vhdl:225:20  */
  assign n1132 = x == 9'b010111101;
  /* fplog32.vhdl:226:20  */
  assign n1135 = x == 9'b010111110;
  /* fplog32.vhdl:227:20  */
  assign n1138 = x == 9'b010111111;
  /* fplog32.vhdl:228:20  */
  assign n1141 = x == 9'b011000000;
  /* fplog32.vhdl:229:20  */
  assign n1144 = x == 9'b011000001;
  /* fplog32.vhdl:230:20  */
  assign n1147 = x == 9'b011000010;
  /* fplog32.vhdl:231:20  */
  assign n1150 = x == 9'b011000011;
  /* fplog32.vhdl:232:20  */
  assign n1153 = x == 9'b011000100;
  /* fplog32.vhdl:233:20  */
  assign n1156 = x == 9'b011000101;
  /* fplog32.vhdl:234:20  */
  assign n1159 = x == 9'b011000110;
  /* fplog32.vhdl:235:20  */
  assign n1162 = x == 9'b011000111;
  /* fplog32.vhdl:236:20  */
  assign n1165 = x == 9'b011001000;
  /* fplog32.vhdl:237:20  */
  assign n1168 = x == 9'b011001001;
  /* fplog32.vhdl:238:20  */
  assign n1171 = x == 9'b011001010;
  /* fplog32.vhdl:239:20  */
  assign n1174 = x == 9'b011001011;
  /* fplog32.vhdl:240:20  */
  assign n1177 = x == 9'b011001100;
  /* fplog32.vhdl:241:20  */
  assign n1180 = x == 9'b011001101;
  /* fplog32.vhdl:242:20  */
  assign n1183 = x == 9'b011001110;
  /* fplog32.vhdl:243:20  */
  assign n1186 = x == 9'b011001111;
  /* fplog32.vhdl:244:20  */
  assign n1189 = x == 9'b011010000;
  /* fplog32.vhdl:245:20  */
  assign n1192 = x == 9'b011010001;
  /* fplog32.vhdl:246:20  */
  assign n1195 = x == 9'b011010010;
  /* fplog32.vhdl:247:20  */
  assign n1198 = x == 9'b011010011;
  /* fplog32.vhdl:248:20  */
  assign n1201 = x == 9'b011010100;
  /* fplog32.vhdl:249:20  */
  assign n1204 = x == 9'b011010101;
  /* fplog32.vhdl:250:20  */
  assign n1207 = x == 9'b011010110;
  /* fplog32.vhdl:251:20  */
  assign n1210 = x == 9'b011010111;
  /* fplog32.vhdl:252:20  */
  assign n1213 = x == 9'b011011000;
  /* fplog32.vhdl:253:20  */
  assign n1216 = x == 9'b011011001;
  /* fplog32.vhdl:254:20  */
  assign n1219 = x == 9'b011011010;
  /* fplog32.vhdl:255:20  */
  assign n1222 = x == 9'b011011011;
  /* fplog32.vhdl:256:20  */
  assign n1225 = x == 9'b011011100;
  /* fplog32.vhdl:257:20  */
  assign n1228 = x == 9'b011011101;
  /* fplog32.vhdl:258:20  */
  assign n1231 = x == 9'b011011110;
  /* fplog32.vhdl:259:20  */
  assign n1234 = x == 9'b011011111;
  /* fplog32.vhdl:260:20  */
  assign n1237 = x == 9'b011100000;
  /* fplog32.vhdl:261:20  */
  assign n1240 = x == 9'b011100001;
  /* fplog32.vhdl:262:20  */
  assign n1243 = x == 9'b011100010;
  /* fplog32.vhdl:263:20  */
  assign n1246 = x == 9'b011100011;
  /* fplog32.vhdl:264:20  */
  assign n1249 = x == 9'b011100100;
  /* fplog32.vhdl:265:20  */
  assign n1252 = x == 9'b011100101;
  /* fplog32.vhdl:266:20  */
  assign n1255 = x == 9'b011100110;
  /* fplog32.vhdl:267:20  */
  assign n1258 = x == 9'b011100111;
  /* fplog32.vhdl:268:20  */
  assign n1261 = x == 9'b011101000;
  /* fplog32.vhdl:269:20  */
  assign n1264 = x == 9'b011101001;
  /* fplog32.vhdl:270:20  */
  assign n1267 = x == 9'b011101010;
  /* fplog32.vhdl:271:20  */
  assign n1270 = x == 9'b011101011;
  /* fplog32.vhdl:272:20  */
  assign n1273 = x == 9'b011101100;
  /* fplog32.vhdl:273:20  */
  assign n1276 = x == 9'b011101101;
  /* fplog32.vhdl:274:20  */
  assign n1279 = x == 9'b011101110;
  /* fplog32.vhdl:275:20  */
  assign n1282 = x == 9'b011101111;
  /* fplog32.vhdl:276:20  */
  assign n1285 = x == 9'b011110000;
  /* fplog32.vhdl:277:20  */
  assign n1288 = x == 9'b011110001;
  /* fplog32.vhdl:278:20  */
  assign n1291 = x == 9'b011110010;
  /* fplog32.vhdl:279:20  */
  assign n1294 = x == 9'b011110011;
  /* fplog32.vhdl:280:20  */
  assign n1297 = x == 9'b011110100;
  /* fplog32.vhdl:281:20  */
  assign n1300 = x == 9'b011110101;
  /* fplog32.vhdl:282:20  */
  assign n1303 = x == 9'b011110110;
  /* fplog32.vhdl:283:20  */
  assign n1306 = x == 9'b011110111;
  /* fplog32.vhdl:284:20  */
  assign n1309 = x == 9'b011111000;
  /* fplog32.vhdl:285:20  */
  assign n1312 = x == 9'b011111001;
  /* fplog32.vhdl:286:20  */
  assign n1315 = x == 9'b011111010;
  /* fplog32.vhdl:287:20  */
  assign n1318 = x == 9'b011111011;
  /* fplog32.vhdl:288:20  */
  assign n1321 = x == 9'b011111100;
  /* fplog32.vhdl:289:20  */
  assign n1324 = x == 9'b011111101;
  /* fplog32.vhdl:290:20  */
  assign n1327 = x == 9'b011111110;
  /* fplog32.vhdl:291:20  */
  assign n1330 = x == 9'b011111111;
  /* fplog32.vhdl:292:20  */
  assign n1333 = x == 9'b100000000;
  /* fplog32.vhdl:293:20  */
  assign n1336 = x == 9'b100000001;
  /* fplog32.vhdl:294:20  */
  assign n1339 = x == 9'b100000010;
  /* fplog32.vhdl:295:20  */
  assign n1342 = x == 9'b100000011;
  /* fplog32.vhdl:296:20  */
  assign n1345 = x == 9'b100000100;
  /* fplog32.vhdl:297:20  */
  assign n1348 = x == 9'b100000101;
  /* fplog32.vhdl:298:20  */
  assign n1351 = x == 9'b100000110;
  /* fplog32.vhdl:299:20  */
  assign n1354 = x == 9'b100000111;
  /* fplog32.vhdl:300:20  */
  assign n1357 = x == 9'b100001000;
  /* fplog32.vhdl:301:20  */
  assign n1360 = x == 9'b100001001;
  /* fplog32.vhdl:302:20  */
  assign n1363 = x == 9'b100001010;
  /* fplog32.vhdl:303:20  */
  assign n1366 = x == 9'b100001011;
  /* fplog32.vhdl:304:20  */
  assign n1369 = x == 9'b100001100;
  /* fplog32.vhdl:305:20  */
  assign n1372 = x == 9'b100001101;
  /* fplog32.vhdl:306:20  */
  assign n1375 = x == 9'b100001110;
  /* fplog32.vhdl:307:20  */
  assign n1378 = x == 9'b100001111;
  /* fplog32.vhdl:308:20  */
  assign n1381 = x == 9'b100010000;
  /* fplog32.vhdl:309:20  */
  assign n1384 = x == 9'b100010001;
  /* fplog32.vhdl:310:20  */
  assign n1387 = x == 9'b100010010;
  /* fplog32.vhdl:311:20  */
  assign n1390 = x == 9'b100010011;
  /* fplog32.vhdl:312:20  */
  assign n1393 = x == 9'b100010100;
  /* fplog32.vhdl:313:20  */
  assign n1396 = x == 9'b100010101;
  /* fplog32.vhdl:314:20  */
  assign n1399 = x == 9'b100010110;
  /* fplog32.vhdl:315:20  */
  assign n1402 = x == 9'b100010111;
  /* fplog32.vhdl:316:20  */
  assign n1405 = x == 9'b100011000;
  /* fplog32.vhdl:317:20  */
  assign n1408 = x == 9'b100011001;
  /* fplog32.vhdl:318:20  */
  assign n1411 = x == 9'b100011010;
  /* fplog32.vhdl:319:20  */
  assign n1414 = x == 9'b100011011;
  /* fplog32.vhdl:320:20  */
  assign n1417 = x == 9'b100011100;
  /* fplog32.vhdl:321:20  */
  assign n1420 = x == 9'b100011101;
  /* fplog32.vhdl:322:20  */
  assign n1423 = x == 9'b100011110;
  /* fplog32.vhdl:323:20  */
  assign n1426 = x == 9'b100011111;
  /* fplog32.vhdl:324:20  */
  assign n1429 = x == 9'b100100000;
  /* fplog32.vhdl:325:20  */
  assign n1432 = x == 9'b100100001;
  /* fplog32.vhdl:326:20  */
  assign n1435 = x == 9'b100100010;
  /* fplog32.vhdl:327:20  */
  assign n1438 = x == 9'b100100011;
  /* fplog32.vhdl:328:20  */
  assign n1441 = x == 9'b100100100;
  /* fplog32.vhdl:329:20  */
  assign n1444 = x == 9'b100100101;
  /* fplog32.vhdl:330:20  */
  assign n1447 = x == 9'b100100110;
  /* fplog32.vhdl:331:20  */
  assign n1450 = x == 9'b100100111;
  /* fplog32.vhdl:332:20  */
  assign n1453 = x == 9'b100101000;
  /* fplog32.vhdl:333:20  */
  assign n1456 = x == 9'b100101001;
  /* fplog32.vhdl:334:20  */
  assign n1459 = x == 9'b100101010;
  /* fplog32.vhdl:335:20  */
  assign n1462 = x == 9'b100101011;
  /* fplog32.vhdl:336:20  */
  assign n1465 = x == 9'b100101100;
  /* fplog32.vhdl:337:20  */
  assign n1468 = x == 9'b100101101;
  /* fplog32.vhdl:338:20  */
  assign n1471 = x == 9'b100101110;
  /* fplog32.vhdl:339:20  */
  assign n1474 = x == 9'b100101111;
  /* fplog32.vhdl:340:20  */
  assign n1477 = x == 9'b100110000;
  /* fplog32.vhdl:341:20  */
  assign n1480 = x == 9'b100110001;
  /* fplog32.vhdl:342:20  */
  assign n1483 = x == 9'b100110010;
  /* fplog32.vhdl:343:20  */
  assign n1486 = x == 9'b100110011;
  /* fplog32.vhdl:344:20  */
  assign n1489 = x == 9'b100110100;
  /* fplog32.vhdl:345:20  */
  assign n1492 = x == 9'b100110101;
  /* fplog32.vhdl:346:20  */
  assign n1495 = x == 9'b100110110;
  /* fplog32.vhdl:347:20  */
  assign n1498 = x == 9'b100110111;
  /* fplog32.vhdl:348:20  */
  assign n1501 = x == 9'b100111000;
  /* fplog32.vhdl:349:20  */
  assign n1504 = x == 9'b100111001;
  /* fplog32.vhdl:350:20  */
  assign n1507 = x == 9'b100111010;
  /* fplog32.vhdl:351:20  */
  assign n1510 = x == 9'b100111011;
  /* fplog32.vhdl:352:20  */
  assign n1513 = x == 9'b100111100;
  /* fplog32.vhdl:353:20  */
  assign n1516 = x == 9'b100111101;
  /* fplog32.vhdl:354:20  */
  assign n1519 = x == 9'b100111110;
  /* fplog32.vhdl:355:20  */
  assign n1522 = x == 9'b100111111;
  /* fplog32.vhdl:356:20  */
  assign n1525 = x == 9'b101000000;
  /* fplog32.vhdl:357:20  */
  assign n1528 = x == 9'b101000001;
  /* fplog32.vhdl:358:20  */
  assign n1531 = x == 9'b101000010;
  /* fplog32.vhdl:359:20  */
  assign n1534 = x == 9'b101000011;
  /* fplog32.vhdl:360:20  */
  assign n1537 = x == 9'b101000100;
  /* fplog32.vhdl:361:20  */
  assign n1540 = x == 9'b101000101;
  /* fplog32.vhdl:362:20  */
  assign n1543 = x == 9'b101000110;
  /* fplog32.vhdl:363:20  */
  assign n1546 = x == 9'b101000111;
  /* fplog32.vhdl:364:20  */
  assign n1549 = x == 9'b101001000;
  /* fplog32.vhdl:365:20  */
  assign n1552 = x == 9'b101001001;
  /* fplog32.vhdl:366:20  */
  assign n1555 = x == 9'b101001010;
  /* fplog32.vhdl:367:20  */
  assign n1558 = x == 9'b101001011;
  /* fplog32.vhdl:368:20  */
  assign n1561 = x == 9'b101001100;
  /* fplog32.vhdl:369:20  */
  assign n1564 = x == 9'b101001101;
  /* fplog32.vhdl:370:20  */
  assign n1567 = x == 9'b101001110;
  /* fplog32.vhdl:371:20  */
  assign n1570 = x == 9'b101001111;
  /* fplog32.vhdl:372:20  */
  assign n1573 = x == 9'b101010000;
  /* fplog32.vhdl:373:20  */
  assign n1576 = x == 9'b101010001;
  /* fplog32.vhdl:374:20  */
  assign n1579 = x == 9'b101010010;
  /* fplog32.vhdl:375:20  */
  assign n1582 = x == 9'b101010011;
  /* fplog32.vhdl:376:20  */
  assign n1585 = x == 9'b101010100;
  /* fplog32.vhdl:377:20  */
  assign n1588 = x == 9'b101010101;
  /* fplog32.vhdl:378:20  */
  assign n1591 = x == 9'b101010110;
  /* fplog32.vhdl:379:20  */
  assign n1594 = x == 9'b101010111;
  /* fplog32.vhdl:380:20  */
  assign n1597 = x == 9'b101011000;
  /* fplog32.vhdl:381:20  */
  assign n1600 = x == 9'b101011001;
  /* fplog32.vhdl:382:20  */
  assign n1603 = x == 9'b101011010;
  /* fplog32.vhdl:383:20  */
  assign n1606 = x == 9'b101011011;
  /* fplog32.vhdl:384:20  */
  assign n1609 = x == 9'b101011100;
  /* fplog32.vhdl:385:20  */
  assign n1612 = x == 9'b101011101;
  /* fplog32.vhdl:386:20  */
  assign n1615 = x == 9'b101011110;
  /* fplog32.vhdl:387:20  */
  assign n1618 = x == 9'b101011111;
  /* fplog32.vhdl:388:20  */
  assign n1621 = x == 9'b101100000;
  /* fplog32.vhdl:389:20  */
  assign n1624 = x == 9'b101100001;
  /* fplog32.vhdl:390:20  */
  assign n1627 = x == 9'b101100010;
  /* fplog32.vhdl:391:20  */
  assign n1630 = x == 9'b101100011;
  /* fplog32.vhdl:392:20  */
  assign n1633 = x == 9'b101100100;
  /* fplog32.vhdl:393:20  */
  assign n1636 = x == 9'b101100101;
  /* fplog32.vhdl:394:20  */
  assign n1639 = x == 9'b101100110;
  /* fplog32.vhdl:395:20  */
  assign n1642 = x == 9'b101100111;
  /* fplog32.vhdl:396:20  */
  assign n1645 = x == 9'b101101000;
  /* fplog32.vhdl:397:20  */
  assign n1648 = x == 9'b101101001;
  /* fplog32.vhdl:398:20  */
  assign n1651 = x == 9'b101101010;
  /* fplog32.vhdl:399:20  */
  assign n1654 = x == 9'b101101011;
  /* fplog32.vhdl:400:20  */
  assign n1657 = x == 9'b101101100;
  /* fplog32.vhdl:401:20  */
  assign n1660 = x == 9'b101101101;
  /* fplog32.vhdl:402:20  */
  assign n1663 = x == 9'b101101110;
  /* fplog32.vhdl:403:20  */
  assign n1666 = x == 9'b101101111;
  /* fplog32.vhdl:404:20  */
  assign n1669 = x == 9'b101110000;
  /* fplog32.vhdl:405:20  */
  assign n1672 = x == 9'b101110001;
  /* fplog32.vhdl:406:20  */
  assign n1675 = x == 9'b101110010;
  /* fplog32.vhdl:407:20  */
  assign n1678 = x == 9'b101110011;
  /* fplog32.vhdl:408:20  */
  assign n1681 = x == 9'b101110100;
  /* fplog32.vhdl:409:20  */
  assign n1684 = x == 9'b101110101;
  /* fplog32.vhdl:410:20  */
  assign n1687 = x == 9'b101110110;
  /* fplog32.vhdl:411:20  */
  assign n1690 = x == 9'b101110111;
  /* fplog32.vhdl:412:20  */
  assign n1693 = x == 9'b101111000;
  /* fplog32.vhdl:413:20  */
  assign n1696 = x == 9'b101111001;
  /* fplog32.vhdl:414:20  */
  assign n1699 = x == 9'b101111010;
  /* fplog32.vhdl:415:20  */
  assign n1702 = x == 9'b101111011;
  /* fplog32.vhdl:416:20  */
  assign n1705 = x == 9'b101111100;
  /* fplog32.vhdl:417:20  */
  assign n1708 = x == 9'b101111101;
  /* fplog32.vhdl:418:20  */
  assign n1711 = x == 9'b101111110;
  /* fplog32.vhdl:419:20  */
  assign n1714 = x == 9'b101111111;
  /* fplog32.vhdl:420:20  */
  assign n1717 = x == 9'b110000000;
  /* fplog32.vhdl:421:20  */
  assign n1720 = x == 9'b110000001;
  /* fplog32.vhdl:422:20  */
  assign n1723 = x == 9'b110000010;
  /* fplog32.vhdl:423:20  */
  assign n1726 = x == 9'b110000011;
  /* fplog32.vhdl:424:20  */
  assign n1729 = x == 9'b110000100;
  /* fplog32.vhdl:425:20  */
  assign n1732 = x == 9'b110000101;
  /* fplog32.vhdl:426:20  */
  assign n1735 = x == 9'b110000110;
  /* fplog32.vhdl:427:20  */
  assign n1738 = x == 9'b110000111;
  /* fplog32.vhdl:428:20  */
  assign n1741 = x == 9'b110001000;
  /* fplog32.vhdl:429:20  */
  assign n1744 = x == 9'b110001001;
  /* fplog32.vhdl:430:20  */
  assign n1747 = x == 9'b110001010;
  /* fplog32.vhdl:431:20  */
  assign n1750 = x == 9'b110001011;
  /* fplog32.vhdl:432:20  */
  assign n1753 = x == 9'b110001100;
  /* fplog32.vhdl:433:20  */
  assign n1756 = x == 9'b110001101;
  /* fplog32.vhdl:434:20  */
  assign n1759 = x == 9'b110001110;
  /* fplog32.vhdl:435:20  */
  assign n1762 = x == 9'b110001111;
  /* fplog32.vhdl:436:20  */
  assign n1765 = x == 9'b110010000;
  /* fplog32.vhdl:437:20  */
  assign n1768 = x == 9'b110010001;
  /* fplog32.vhdl:438:20  */
  assign n1771 = x == 9'b110010010;
  /* fplog32.vhdl:439:20  */
  assign n1774 = x == 9'b110010011;
  /* fplog32.vhdl:440:20  */
  assign n1777 = x == 9'b110010100;
  /* fplog32.vhdl:441:20  */
  assign n1780 = x == 9'b110010101;
  /* fplog32.vhdl:442:20  */
  assign n1783 = x == 9'b110010110;
  /* fplog32.vhdl:443:20  */
  assign n1786 = x == 9'b110010111;
  /* fplog32.vhdl:444:20  */
  assign n1789 = x == 9'b110011000;
  /* fplog32.vhdl:445:20  */
  assign n1792 = x == 9'b110011001;
  /* fplog32.vhdl:446:20  */
  assign n1795 = x == 9'b110011010;
  /* fplog32.vhdl:447:20  */
  assign n1798 = x == 9'b110011011;
  /* fplog32.vhdl:448:20  */
  assign n1801 = x == 9'b110011100;
  /* fplog32.vhdl:449:20  */
  assign n1804 = x == 9'b110011101;
  /* fplog32.vhdl:450:20  */
  assign n1807 = x == 9'b110011110;
  /* fplog32.vhdl:451:20  */
  assign n1810 = x == 9'b110011111;
  /* fplog32.vhdl:452:20  */
  assign n1813 = x == 9'b110100000;
  /* fplog32.vhdl:453:20  */
  assign n1816 = x == 9'b110100001;
  /* fplog32.vhdl:454:20  */
  assign n1819 = x == 9'b110100010;
  /* fplog32.vhdl:455:20  */
  assign n1822 = x == 9'b110100011;
  /* fplog32.vhdl:456:20  */
  assign n1825 = x == 9'b110100100;
  /* fplog32.vhdl:457:20  */
  assign n1828 = x == 9'b110100101;
  /* fplog32.vhdl:458:20  */
  assign n1831 = x == 9'b110100110;
  /* fplog32.vhdl:459:20  */
  assign n1834 = x == 9'b110100111;
  /* fplog32.vhdl:460:20  */
  assign n1837 = x == 9'b110101000;
  /* fplog32.vhdl:461:20  */
  assign n1840 = x == 9'b110101001;
  /* fplog32.vhdl:462:20  */
  assign n1843 = x == 9'b110101010;
  /* fplog32.vhdl:463:20  */
  assign n1846 = x == 9'b110101011;
  /* fplog32.vhdl:464:20  */
  assign n1849 = x == 9'b110101100;
  /* fplog32.vhdl:465:20  */
  assign n1852 = x == 9'b110101101;
  /* fplog32.vhdl:466:20  */
  assign n1855 = x == 9'b110101110;
  /* fplog32.vhdl:467:20  */
  assign n1858 = x == 9'b110101111;
  /* fplog32.vhdl:468:20  */
  assign n1861 = x == 9'b110110000;
  /* fplog32.vhdl:469:20  */
  assign n1864 = x == 9'b110110001;
  /* fplog32.vhdl:470:20  */
  assign n1867 = x == 9'b110110010;
  /* fplog32.vhdl:471:20  */
  assign n1870 = x == 9'b110110011;
  /* fplog32.vhdl:472:20  */
  assign n1873 = x == 9'b110110100;
  /* fplog32.vhdl:473:20  */
  assign n1876 = x == 9'b110110101;
  /* fplog32.vhdl:474:20  */
  assign n1879 = x == 9'b110110110;
  /* fplog32.vhdl:475:20  */
  assign n1882 = x == 9'b110110111;
  /* fplog32.vhdl:476:20  */
  assign n1885 = x == 9'b110111000;
  /* fplog32.vhdl:477:20  */
  assign n1888 = x == 9'b110111001;
  /* fplog32.vhdl:478:20  */
  assign n1891 = x == 9'b110111010;
  /* fplog32.vhdl:479:20  */
  assign n1894 = x == 9'b110111011;
  /* fplog32.vhdl:480:20  */
  assign n1897 = x == 9'b110111100;
  /* fplog32.vhdl:481:20  */
  assign n1900 = x == 9'b110111101;
  /* fplog32.vhdl:482:20  */
  assign n1903 = x == 9'b110111110;
  /* fplog32.vhdl:483:20  */
  assign n1906 = x == 9'b110111111;
  /* fplog32.vhdl:484:20  */
  assign n1909 = x == 9'b111000000;
  /* fplog32.vhdl:485:20  */
  assign n1912 = x == 9'b111000001;
  /* fplog32.vhdl:486:20  */
  assign n1915 = x == 9'b111000010;
  /* fplog32.vhdl:487:20  */
  assign n1918 = x == 9'b111000011;
  /* fplog32.vhdl:488:20  */
  assign n1921 = x == 9'b111000100;
  /* fplog32.vhdl:489:20  */
  assign n1924 = x == 9'b111000101;
  /* fplog32.vhdl:490:20  */
  assign n1927 = x == 9'b111000110;
  /* fplog32.vhdl:491:20  */
  assign n1930 = x == 9'b111000111;
  /* fplog32.vhdl:492:20  */
  assign n1933 = x == 9'b111001000;
  /* fplog32.vhdl:493:20  */
  assign n1936 = x == 9'b111001001;
  /* fplog32.vhdl:494:20  */
  assign n1939 = x == 9'b111001010;
  /* fplog32.vhdl:495:20  */
  assign n1942 = x == 9'b111001011;
  /* fplog32.vhdl:496:20  */
  assign n1945 = x == 9'b111001100;
  /* fplog32.vhdl:497:20  */
  assign n1948 = x == 9'b111001101;
  /* fplog32.vhdl:498:20  */
  assign n1951 = x == 9'b111001110;
  /* fplog32.vhdl:499:20  */
  assign n1954 = x == 9'b111001111;
  /* fplog32.vhdl:500:20  */
  assign n1957 = x == 9'b111010000;
  /* fplog32.vhdl:501:20  */
  assign n1960 = x == 9'b111010001;
  /* fplog32.vhdl:502:20  */
  assign n1963 = x == 9'b111010010;
  /* fplog32.vhdl:503:20  */
  assign n1966 = x == 9'b111010011;
  /* fplog32.vhdl:504:20  */
  assign n1969 = x == 9'b111010100;
  /* fplog32.vhdl:505:20  */
  assign n1972 = x == 9'b111010101;
  /* fplog32.vhdl:506:20  */
  assign n1975 = x == 9'b111010110;
  /* fplog32.vhdl:507:20  */
  assign n1978 = x == 9'b111010111;
  /* fplog32.vhdl:508:20  */
  assign n1981 = x == 9'b111011000;
  /* fplog32.vhdl:509:20  */
  assign n1984 = x == 9'b111011001;
  /* fplog32.vhdl:510:20  */
  assign n1987 = x == 9'b111011010;
  /* fplog32.vhdl:511:20  */
  assign n1990 = x == 9'b111011011;
  /* fplog32.vhdl:512:20  */
  assign n1993 = x == 9'b111011100;
  /* fplog32.vhdl:513:20  */
  assign n1996 = x == 9'b111011101;
  /* fplog32.vhdl:514:20  */
  assign n1999 = x == 9'b111011110;
  /* fplog32.vhdl:515:20  */
  assign n2002 = x == 9'b111011111;
  /* fplog32.vhdl:516:20  */
  assign n2005 = x == 9'b111100000;
  /* fplog32.vhdl:517:20  */
  assign n2008 = x == 9'b111100001;
  /* fplog32.vhdl:518:20  */
  assign n2011 = x == 9'b111100010;
  /* fplog32.vhdl:519:20  */
  assign n2014 = x == 9'b111100011;
  /* fplog32.vhdl:520:20  */
  assign n2017 = x == 9'b111100100;
  /* fplog32.vhdl:521:20  */
  assign n2020 = x == 9'b111100101;
  /* fplog32.vhdl:522:20  */
  assign n2023 = x == 9'b111100110;
  /* fplog32.vhdl:523:20  */
  assign n2026 = x == 9'b111100111;
  /* fplog32.vhdl:524:20  */
  assign n2029 = x == 9'b111101000;
  /* fplog32.vhdl:525:20  */
  assign n2032 = x == 9'b111101001;
  /* fplog32.vhdl:526:20  */
  assign n2035 = x == 9'b111101010;
  /* fplog32.vhdl:527:20  */
  assign n2038 = x == 9'b111101011;
  /* fplog32.vhdl:528:20  */
  assign n2041 = x == 9'b111101100;
  /* fplog32.vhdl:529:20  */
  assign n2044 = x == 9'b111101101;
  /* fplog32.vhdl:530:20  */
  assign n2047 = x == 9'b111101110;
  /* fplog32.vhdl:531:20  */
  assign n2050 = x == 9'b111101111;
  /* fplog32.vhdl:532:20  */
  assign n2053 = x == 9'b111110000;
  /* fplog32.vhdl:533:20  */
  assign n2056 = x == 9'b111110001;
  /* fplog32.vhdl:534:20  */
  assign n2059 = x == 9'b111110010;
  /* fplog32.vhdl:535:20  */
  assign n2062 = x == 9'b111110011;
  /* fplog32.vhdl:536:20  */
  assign n2065 = x == 9'b111110100;
  /* fplog32.vhdl:537:20  */
  assign n2068 = x == 9'b111110101;
  /* fplog32.vhdl:538:20  */
  assign n2071 = x == 9'b111110110;
  /* fplog32.vhdl:539:20  */
  assign n2074 = x == 9'b111110111;
  /* fplog32.vhdl:540:20  */
  assign n2077 = x == 9'b111111000;
  /* fplog32.vhdl:541:20  */
  assign n2080 = x == 9'b111111001;
  /* fplog32.vhdl:542:20  */
  assign n2083 = x == 9'b111111010;
  /* fplog32.vhdl:543:20  */
  assign n2086 = x == 9'b111111011;
  /* fplog32.vhdl:544:20  */
  assign n2089 = x == 9'b111111100;
  /* fplog32.vhdl:545:20  */
  assign n2092 = x == 9'b111111101;
  /* fplog32.vhdl:546:20  */
  assign n2095 = x == 9'b111111110;
  /* fplog32.vhdl:547:20  */
  assign n2098 = x == 9'b111111111;
  assign n2100 = {n2098, n2095, n2092, n2089, n2086, n2083, n2080, n2077, n2074, n2071, n2068, n2065, n2062, n2059, n2056, n2053, n2050, n2047, n2044, n2041, n2038, n2035, n2032, n2029, n2026, n2023, n2020, n2017, n2014, n2011, n2008, n2005, n2002, n1999, n1996, n1993, n1990, n1987, n1984, n1981, n1978, n1975, n1972, n1969, n1966, n1963, n1960, n1957, n1954, n1951, n1948, n1945, n1942, n1939, n1936, n1933, n1930, n1927, n1924, n1921, n1918, n1915, n1912, n1909, n1906, n1903, n1900, n1897, n1894, n1891, n1888, n1885, n1882, n1879, n1876, n1873, n1870, n1867, n1864, n1861, n1858, n1855, n1852, n1849, n1846, n1843, n1840, n1837, n1834, n1831, n1828, n1825, n1822, n1819, n1816, n1813, n1810, n1807, n1804, n1801, n1798, n1795, n1792, n1789, n1786, n1783, n1780, n1777, n1774, n1771, n1768, n1765, n1762, n1759, n1756, n1753, n1750, n1747, n1744, n1741, n1738, n1735, n1732, n1729, n1726, n1723, n1720, n1717, n1714, n1711, n1708, n1705, n1702, n1699, n1696, n1693, n1690, n1687, n1684, n1681, n1678, n1675, n1672, n1669, n1666, n1663, n1660, n1657, n1654, n1651, n1648, n1645, n1642, n1639, n1636, n1633, n1630, n1627, n1624, n1621, n1618, n1615, n1612, n1609, n1606, n1603, n1600, n1597, n1594, n1591, n1588, n1585, n1582, n1579, n1576, n1573, n1570, n1567, n1564, n1561, n1558, n1555, n1552, n1549, n1546, n1543, n1540, n1537, n1534, n1531, n1528, n1525, n1522, n1519, n1516, n1513, n1510, n1507, n1504, n1501, n1498, n1495, n1492, n1489, n1486, n1483, n1480, n1477, n1474, n1471, n1468, n1465, n1462, n1459, n1456, n1453, n1450, n1447, n1444, n1441, n1438, n1435, n1432, n1429, n1426, n1423, n1420, n1417, n1414, n1411, n1408, n1405, n1402, n1399, n1396, n1393, n1390, n1387, n1384, n1381, n1378, n1375, n1372, n1369, n1366, n1363, n1360, n1357, n1354, n1351, n1348, n1345, n1342, n1339, n1336, n1333, n1330, n1327, n1324, n1321, n1318, n1315, n1312, n1309, n1306, n1303, n1300, n1297, n1294, n1291, n1288, n1285, n1282, n1279, n1276, n1273, n1270, n1267, n1264, n1261, n1258, n1255, n1252, n1249, n1246, n1243, n1240, n1237, n1234, n1231, n1228, n1225, n1222, n1219, n1216, n1213, n1210, n1207, n1204, n1201, n1198, n1195, n1192, n1189, n1186, n1183, n1180, n1177, n1174, n1171, n1168, n1165, n1162, n1159, n1156, n1153, n1150, n1147, n1144, n1141, n1138, n1135, n1132, n1129, n1126, n1123, n1120, n1117, n1114, n1111, n1108, n1105, n1102, n1099, n1096, n1093, n1090, n1087, n1084, n1081, n1078, n1075, n1072, n1069, n1066, n1063, n1060, n1057, n1054, n1051, n1048, n1045, n1042, n1039, n1036, n1033, n1030, n1027, n1024, n1021, n1018, n1015, n1012, n1009, n1006, n1003, n1000, n997, n994, n991, n988, n985, n982, n979, n976, n973, n970, n967, n964, n961, n958, n955, n952, n949, n946, n943, n940, n937, n934, n931, n928, n925, n922, n919, n916, n913, n910, n907, n904, n901, n898, n895, n892, n889, n886, n883, n880, n877, n874, n871, n868, n865, n862, n859, n856, n853, n850, n847, n844, n841, n838, n835, n832, n829, n826, n823, n820, n817, n814, n811, n808, n805, n802, n799, n796, n793, n790, n787, n784, n781, n778, n775, n772, n769, n766, n763, n760, n757, n754, n751, n748, n745, n742, n739, n736, n733, n730, n727, n724, n721, n718, n715, n712, n709, n706, n703, n700, n697, n694, n691, n688, n685, n682, n679, n676, n673, n670, n667, n664, n661, n658, n655, n652, n649, n646, n643, n640, n637, n634, n631, n628, n625, n622, n619, n616, n613, n610, n607, n604, n601, n598, n595, n592, n589, n586, n583, n580, n577, n574, n571, n568, n565};
  /* fplog32.vhdl:35:4  */
  always @*
    case (n2100)
      512'b10000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b1000000001;
      512'b01000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b1000000010;
      512'b00100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b1000000010;
      512'b00010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b1000000011;
      512'b00001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b1000000011;
      512'b00000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b1000000100;
      512'b00000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b1000000100;
      512'b00000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b1000000101;
      512'b00000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b1000000101;
      512'b00000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b1000000110;
      512'b00000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b1000000110;
      512'b00000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b1000000111;
      512'b00000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b1000000111;
      512'b00000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b1000001000;
      512'b00000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b1000001000;
      512'b00000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b1000001001;
      512'b00000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b1000001001;
      512'b00000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b1000001010;
      512'b00000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b1000001010;
      512'b00000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b1000001011;
      512'b00000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b1000001011;
      512'b00000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b1000001100;
      512'b00000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b1000001100;
      512'b00000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b1000001101;
      512'b00000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b1000001101;
      512'b00000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b1000001110;
      512'b00000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b1000001110;
      512'b00000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b1000001111;
      512'b00000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b1000001111;
      512'b00000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b1000010000;
      512'b00000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b1000010000;
      512'b00000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b1000010001;
      512'b00000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b1000010010;
      512'b00000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b1000010010;
      512'b00000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b1000010011;
      512'b00000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b1000010011;
      512'b00000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b1000010100;
      512'b00000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b1000010100;
      512'b00000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b1000010101;
      512'b00000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b1000010101;
      512'b00000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b1000010110;
      512'b00000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b1000010110;
      512'b00000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b1000010111;
      512'b00000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b1000010111;
      512'b00000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b1000011000;
      512'b00000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b1000011001;
      512'b00000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b1000011001;
      512'b00000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b1000011010;
      512'b00000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b1000011010;
      512'b00000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b1000011011;
      512'b00000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b1000011011;
      512'b00000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b1000011100;
      512'b00000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b1000011100;
      512'b00000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b1000011101;
      512'b00000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b1000011110;
      512'b00000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b1000011110;
      512'b00000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b1000011111;
      512'b00000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b1000011111;
      512'b00000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b1000100000;
      512'b00000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b1000100000;
      512'b00000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b1000100001;
      512'b00000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b1000100001;
      512'b00000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b1000100010;
      512'b00000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b1000100011;
      512'b00000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b1000100011;
      512'b00000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b1000100100;
      512'b00000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b1000100100;
      512'b00000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b1000100101;
      512'b00000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b1000100101;
      512'b00000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b1000100110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b1000100111;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b1000100111;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b1000101000;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b1000101000;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b1000101001;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b1000101010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b1000101010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b1000101011;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b1000101011;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b1000101100;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b1000101100;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b1000101101;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b1000101110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b1000101110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b1000101111;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b1000101111;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b1000110000;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b1000110001;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b1000110001;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b1000110010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b1000110010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b1000110011;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b1000110100;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b1000110100;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b1000110101;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b1000110101;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b1000110110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b1000110111;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b1000110111;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b1000111000;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b1000111001;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b1000111001;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b1000111010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b1000111010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b1000111011;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b1000111100;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b1000111100;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b1000111101;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b1000111101;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b1000111110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b1000111111;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b1000111111;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b1001000000;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b1001000001;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b1001000001;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b1001000010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b1001000011;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b1001000011;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b1001000100;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b1001000100;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b1001000101;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b1001000110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b1001000110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b1001000111;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b1001001000;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b1001001000;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b1001001001;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b1001001010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b1001001010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b1001001011;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b1001001100;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b1001001100;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b1001001101;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b1001001110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b1001001110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b1001001111;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b1001010000;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b1001010000;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b1001010001;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b1001010010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b1001010010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b1001010011;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b1001010100;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b1001010100;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b1001010101;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b1001010110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b1001010110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b1001010111;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b1001011000;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b1001011000;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b1001011001;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b1001011010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b1001011010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b1001011011;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b1001011100;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b1001011101;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b1001011101;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b1001011110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b1001011111;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b1001011111;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b1001100000;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b1001100001;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b1001100001;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b1001100010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b1001100011;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b1001100100;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b1001100100;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b1001100101;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b1001100110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b1001100110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b1001100111;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b1001101000;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b1001101001;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b1001101001;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b1001101010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b1001101011;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b1001101011;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b1001101100;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b1001101101;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b1001101110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b1001101110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b1001101111;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b1001110000;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b1001110001;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b1001110001;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b1001110010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b1001110011;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b1001110100;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b1001110100;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b1001110101;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b1001110110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b1001110111;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b1001110111;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b1001111000;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b1001111001;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b1001111010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b1001111010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b1001111011;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b1001111100;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b1001111101;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b1001111110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b1001111110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b1001111111;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b1010000000;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b1010000001;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b1010000001;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b1010000010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b1010000011;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b1010000100;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b1010000101;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b1010000101;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b1010000110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b1010000111;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b1010001000;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b1010001001;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b1010001001;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b1010001010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b1010001011;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b1010001100;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b1010001101;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b1010001101;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b1010001110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b1010001111;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b1010010000;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b1010010001;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b1010010010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b1010010010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b1010010011;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b1010010100;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b1010010101;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b1010010110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b1010010110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b1010010111;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b1010011000;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b1010011001;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b1010011010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b1010011011;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b1010011100;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b1010011100;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b1010011101;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b1010011110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b1010011111;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b1010100000;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b1010100001;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b1010100010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b1010100010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b1010100011;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b1010100100;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b1010100101;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b1010100110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b1010100111;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b1010101000;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b1010101001;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b1010101001;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b1010101010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b1010101011;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b0101010110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b0101010111;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b0101010111;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b0101011000;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b0101011000;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b0101011001;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b0101011001;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b0101011001;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b0101011010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b0101011010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b0101011011;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b0101011011;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b0101011100;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b0101011100;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b0101011101;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b0101011101;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b0101011110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b0101011110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b0101011110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b0101011111;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b0101011111;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b0101100000;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b0101100000;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b0101100001;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b0101100001;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b0101100010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b0101100010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b0101100011;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b0101100011;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b0101100100;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b0101100100;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b0101100101;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b0101100101;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b0101100110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b0101100110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b0101100111;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b0101100111;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b0101101000;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b0101101000;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b0101101001;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b0101101001;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b0101101010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b0101101010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b0101101011;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b0101101011;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b0101101100;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b0101101100;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b0101101101;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b0101101101;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b0101101110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b0101101110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b0101101111;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b0101101111;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b0101110000;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b0101110000;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b0101110001;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b0101110001;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b0101110010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b0101110010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b0101110011;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b0101110011;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b0101110100;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b0101110100;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b0101110101;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b0101110101;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b0101110110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b0101110110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b0101110111;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b0101111000;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b0101111000;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b0101111001;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b0101111001;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b0101111010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b0101111010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b0101111011;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b0101111011;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b0101111100;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b0101111100;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b0101111101;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b0101111110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b0101111110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b0101111111;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b0101111111;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b0110000000;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b0110000000;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b0110000001;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b0110000001;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b0110000010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b0110000011;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b0110000011;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b0110000100;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b0110000100;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b0110000101;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b0110000101;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b0110000110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b0110000111;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b0110000111;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b0110001000;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b0110001000;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b0110001001;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b0110001010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b0110001010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b0110001011;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b0110001011;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b0110001100;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b0110001100;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b0110001101;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b0110001110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b0110001110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b0110001111;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b0110010000;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b0110010000;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b0110010001;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b0110010001;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b0110010010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b0110010011;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b0110010011;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b0110010100;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b0110010100;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b0110010101;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b0110010110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b0110010110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b0110010111;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b0110011000;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b0110011000;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b0110011001;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b0110011001;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b0110011010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b0110011011;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b0110011011;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b0110011100;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b0110011101;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b0110011101;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b0110011110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b0110011111;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b0110011111;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b0110100000;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b0110100001;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b0110100001;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b0110100010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b0110100011;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b0110100011;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b0110100100;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b0110100101;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b0110100101;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b0110100110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b0110100111;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b0110100111;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b0110101000;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b0110101001;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b0110101001;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b0110101010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b0110101011;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b0110101011;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b0110101100;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b0110101101;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b0110101110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b0110101110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b0110101111;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b0110110000;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b0110110000;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b0110110001;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b0110110010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b0110110011;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b0110110011;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b0110110100;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b0110110101;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b0110110101;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b0110110110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b0110110111;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b0110111000;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b0110111000;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b0110111001;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b0110111010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b0110111011;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b0110111011;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b0110111100;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b0110111101;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b0110111110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b0110111110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b0110111111;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b0111000000;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b0111000001;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b0111000001;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b0111000010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b0111000011;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b0111000100;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b0111000100;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b0111000101;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b0111000110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b0111000111;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b0111001000;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b0111001000;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b0111001001;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b0111001010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000: n2101 = 10'b0111001011;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000: n2101 = 10'b0111001100;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000: n2101 = 10'b0111001100;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000: n2101 = 10'b0111001101;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000: n2101 = 10'b0111001110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000: n2101 = 10'b0111001111;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000: n2101 = 10'b0111010000;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000: n2101 = 10'b0111010000;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000: n2101 = 10'b0111010001;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000: n2101 = 10'b0111010010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000: n2101 = 10'b0111010011;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000: n2101 = 10'b0111010100;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000: n2101 = 10'b0111010101;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000: n2101 = 10'b0111010101;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000: n2101 = 10'b0111010110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000: n2101 = 10'b0111010111;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000: n2101 = 10'b0111011000;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000: n2101 = 10'b0111011001;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000: n2101 = 10'b0111011010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000: n2101 = 10'b0111011011;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000: n2101 = 10'b0111011011;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000: n2101 = 10'b0111011100;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000: n2101 = 10'b0111011101;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000: n2101 = 10'b0111011110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000: n2101 = 10'b0111011111;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000: n2101 = 10'b0111100000;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000: n2101 = 10'b0111100001;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000: n2101 = 10'b0111100001;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000: n2101 = 10'b0111100010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000: n2101 = 10'b0111100011;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000: n2101 = 10'b0111100100;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000: n2101 = 10'b0111100101;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000: n2101 = 10'b0111100110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000: n2101 = 10'b0111100111;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000: n2101 = 10'b0111101000;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000: n2101 = 10'b0111101001;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000: n2101 = 10'b0111101010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000: n2101 = 10'b0111101010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000: n2101 = 10'b0111101011;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000: n2101 = 10'b0111101100;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000: n2101 = 10'b0111101101;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000: n2101 = 10'b0111101110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000: n2101 = 10'b0111101111;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000: n2101 = 10'b0111110000;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000: n2101 = 10'b0111110001;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000: n2101 = 10'b0111110010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000: n2101 = 10'b0111110011;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000: n2101 = 10'b0111110100;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000: n2101 = 10'b0111110101;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000: n2101 = 10'b0111110110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000: n2101 = 10'b0111110111;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000: n2101 = 10'b0111111000;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000: n2101 = 10'b0111111001;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000: n2101 = 10'b0111111010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000: n2101 = 10'b0111111011;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000: n2101 = 10'b0111111100;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000: n2101 = 10'b0111111101;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000: n2101 = 10'b0111111110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100: n2101 = 10'b0111111111;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010: n2101 = 10'b1000000000;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001: n2101 = 10'b1000000000;
      default: n2101 = 10'bX;
    endcase
endmodule

module leftshifter12_by_max_12_freq500_uid6
  (input  clk,
   input  [11:0] x,
   input  [3:0] s,
   output [23:0] r);
  wire [3:0] ps;
  wire [3:0] ps_d1;
  wire [11:0] level0;
  wire [11:0] level0_d1;
  wire [11:0] level0_d2;
  wire [11:0] level0_d3;
  wire [12:0] level1;
  wire [12:0] level1_d1;
  wire [14:0] level2;
  wire [18:0] level3;
  wire [26:0] level4;
  wire [12:0] n533;
  wire n534;
  wire [12:0] n535;
  wire [12:0] n537;
  wire [14:0] n539;
  wire n540;
  wire [14:0] n541;
  wire [14:0] n543;
  wire [18:0] n545;
  wire n546;
  wire [18:0] n547;
  wire [18:0] n549;
  wire [26:0] n551;
  wire n552;
  wire [26:0] n553;
  wire [26:0] n555;
  wire [23:0] n556;
  reg [3:0] n557;
  reg [11:0] n558;
  reg [11:0] n559;
  reg [11:0] n560;
  reg [12:0] n561;
  assign r = n556; //(module output)
  /* fplog32.vhdl:967:12  */
  assign ps_d1 = n557; // (signal)
  /* fplog32.vhdl:969:16  */
  assign level0_d1 = n558; // (signal)
  /* fplog32.vhdl:969:27  */
  assign level0_d2 = n559; // (signal)
  /* fplog32.vhdl:969:38  */
  assign level0_d3 = n560; // (signal)
  /* fplog32.vhdl:971:8  */
  assign level1 = n535; // (signal)
  /* fplog32.vhdl:971:16  */
  assign level1_d1 = n561; // (signal)
  /* fplog32.vhdl:973:8  */
  assign level2 = n541; // (signal)
  /* fplog32.vhdl:975:8  */
  assign level3 = n547; // (signal)
  /* fplog32.vhdl:977:8  */
  assign level4 = n553; // (signal)
  /* fplog32.vhdl:992:23  */
  assign n533 = {level0_d3, 1'b0};
  /* fplog32.vhdl:992:52  */
  assign n534 = ps[0]; // extract
  /* fplog32.vhdl:992:45  */
  assign n535 = n534 ? n533 : n537;
  /* fplog32.vhdl:992:90  */
  assign n537 = {1'b0, level0_d3};
  /* fplog32.vhdl:993:23  */
  assign n539 = {level1_d1, 2'b00};
  /* fplog32.vhdl:993:55  */
  assign n540 = ps_d1[1]; // extract
  /* fplog32.vhdl:993:45  */
  assign n541 = n540 ? n539 : n543;
  /* fplog32.vhdl:993:93  */
  assign n543 = {2'b00, level1_d1};
  /* fplog32.vhdl:994:20  */
  assign n545 = {level2, 4'b0000};
  /* fplog32.vhdl:994:52  */
  assign n546 = ps_d1[2]; // extract
  /* fplog32.vhdl:994:42  */
  assign n547 = n546 ? n545 : n549;
  /* fplog32.vhdl:994:90  */
  assign n549 = {4'b0000, level2};
  /* fplog32.vhdl:995:20  */
  assign n551 = {level3, 8'b00000000};
  /* fplog32.vhdl:995:52  */
  assign n552 = ps_d1[3]; // extract
  /* fplog32.vhdl:995:42  */
  assign n553 = n552 ? n551 : n555;
  /* fplog32.vhdl:995:90  */
  assign n555 = {8'b00000000, level3};
  /* fplog32.vhdl:996:15  */
  assign n556 = level4[23:0]; // extract
  /* fplog32.vhdl:982:10  */
  always @(posedge clk)
    n557 <= ps;
  /* fplog32.vhdl:982:10  */
  always @(posedge clk)
    n558 <= level0;
  /* fplog32.vhdl:982:10  */
  always @(posedge clk)
    n559 <= level0_d1;
  /* fplog32.vhdl:982:10  */
  always @(posedge clk)
    n560 <= level0_d2;
  /* fplog32.vhdl:982:10  */
  always @(posedge clk)
    n561 <= level1;
endmodule

module lzoc_23_freq500_uid4
  (input  clk,
   input  [22:0] i,
   input  ozb,
   output [4:0] o);
  wire sozb;
  wire sozb_d1;
  wire sozb_d2;
  wire [30:0] level5;
  wire [30:0] level5_d1;
  wire digit4;
  wire digit4_d1;
  wire digit4_d2;
  wire [14:0] level4;
  wire [14:0] level4_d1;
  wire digit3;
  wire digit3_d1;
  wire [6:0] level3;
  wire digit2;
  wire [2:0] level2;
  wire [2:0] level2_d1;
  wire [2:0] z;
  wire [1:0] lowbits;
  wire [2:0] outhighbits;
  wire [2:0] outhighbits_d1;
  wire ozb_d1;
  wire ozb_d2;
  wire ozb_d3;
  wire n443;
  wire n444;
  wire n445;
  wire n446;
  wire n447;
  wire n448;
  wire n449;
  wire n450;
  wire [3:0] n451;
  wire [3:0] n452;
  wire [7:0] n453;
  wire [30:0] n454;
  wire [15:0] n456;
  wire [3:0] n457;
  wire [3:0] n458;
  wire [3:0] n459;
  wire [3:0] n460;
  wire [15:0] n461;
  wire n462;
  wire n463;
  wire [14:0] n465;
  wire [14:0] n466;
  wire [14:0] n467;
  wire [7:0] n469;
  wire [3:0] n470;
  wire [3:0] n471;
  wire [7:0] n472;
  wire n473;
  wire n474;
  wire [6:0] n476;
  wire [6:0] n477;
  wire [6:0] n478;
  wire [3:0] n480;
  wire [3:0] n481;
  wire n482;
  wire n483;
  wire [2:0] n485;
  wire [2:0] n486;
  wire [2:0] n487;
  wire n488;
  wire [2:0] n489;
  wire [2:0] n490;
  wire n493;
  wire n496;
  wire n499;
  wire n502;
  wire [3:0] n504;
  reg [1:0] n505;
  wire [1:0] n506;
  wire [2:0] n507;
  wire [4:0] n509;
  reg n510;
  reg n511;
  reg [30:0] n512;
  reg n513;
  reg n514;
  reg [14:0] n515;
  reg n516;
  reg [2:0] n517;
  reg [2:0] n518;
  reg n519;
  reg n520;
  reg n521;
  assign o = n509; //(module output)
  /* fplog32.vhdl:872:8  */
  assign sozb = ozb; // (signal)
  /* fplog32.vhdl:872:14  */
  assign sozb_d1 = n510; // (signal)
  /* fplog32.vhdl:872:23  */
  assign sozb_d2 = n511; // (signal)
  /* fplog32.vhdl:874:8  */
  assign level5 = n454; // (signal)
  /* fplog32.vhdl:874:16  */
  assign level5_d1 = n512; // (signal)
  /* fplog32.vhdl:876:8  */
  assign digit4 = n463; // (signal)
  /* fplog32.vhdl:876:16  */
  assign digit4_d1 = n513; // (signal)
  /* fplog32.vhdl:876:27  */
  assign digit4_d2 = n514; // (signal)
  /* fplog32.vhdl:878:8  */
  assign level4 = n466; // (signal)
  /* fplog32.vhdl:878:16  */
  assign level4_d1 = n515; // (signal)
  /* fplog32.vhdl:880:8  */
  assign digit3 = n474; // (signal)
  /* fplog32.vhdl:880:16  */
  assign digit3_d1 = n516; // (signal)
  /* fplog32.vhdl:882:8  */
  assign level3 = n477; // (signal)
  /* fplog32.vhdl:884:8  */
  assign digit2 = n483; // (signal)
  /* fplog32.vhdl:886:8  */
  assign level2 = n486; // (signal)
  /* fplog32.vhdl:886:16  */
  assign level2_d1 = n517; // (signal)
  /* fplog32.vhdl:888:8  */
  assign z = n489; // (signal)
  /* fplog32.vhdl:890:8  */
  assign lowbits = n505; // (signal)
  /* fplog32.vhdl:892:8  */
  assign outhighbits = n507; // (signal)
  /* fplog32.vhdl:892:21  */
  assign outhighbits_d1 = n518; // (signal)
  /* fplog32.vhdl:894:8  */
  assign ozb_d1 = n519; // (signal)
  /* fplog32.vhdl:894:16  */
  assign ozb_d2 = n520; // (signal)
  /* fplog32.vhdl:894:24  */
  assign ozb_d3 = n521; // (signal)
  /* fplog32.vhdl:916:33  */
  assign n443 = ~sozb;
  /* fplog32.vhdl:916:33  */
  assign n444 = ~sozb;
  /* fplog32.vhdl:916:33  */
  assign n445 = ~sozb;
  /* fplog32.vhdl:916:33  */
  assign n446 = ~sozb;
  /* fplog32.vhdl:916:33  */
  assign n447 = ~sozb;
  /* fplog32.vhdl:916:33  */
  assign n448 = ~sozb;
  /* fplog32.vhdl:916:33  */
  assign n449 = ~sozb;
  /* fplog32.vhdl:916:33  */
  assign n450 = ~sozb;
  assign n451 = {n450, n449, n448, n447};
  assign n452 = {n446, n445, n444, n443};
  assign n453 = {n451, n452};
  /* fplog32.vhdl:916:16  */
  assign n454 = {i, n453};
  /* fplog32.vhdl:918:28  */
  assign n456 = level5[30:15]; // extract
  assign n457 = {sozb, sozb, sozb, sozb};
  assign n458 = {sozb, sozb, sozb, sozb};
  assign n459 = {sozb, sozb, sozb, sozb};
  assign n460 = {sozb, sozb, sozb, sozb};
  assign n461 = {n457, n458, n459, n460};
  /* fplog32.vhdl:918:43  */
  assign n462 = n456 == n461;
  /* fplog32.vhdl:918:17  */
  assign n463 = n462 ? 1'b1 : 1'b0;
  /* fplog32.vhdl:919:22  */
  assign n465 = level5_d1[14:0]; // extract
  /* fplog32.vhdl:919:36  */
  assign n466 = digit4_d1 ? n465 : n467;
  /* fplog32.vhdl:919:69  */
  assign n467 = level5_d1[30:16]; // extract
  /* fplog32.vhdl:920:28  */
  assign n469 = level4[14:7]; // extract
  assign n470 = {sozb_d1, sozb_d1, sozb_d1, sozb_d1};
  assign n471 = {sozb_d1, sozb_d1, sozb_d1, sozb_d1};
  assign n472 = {n470, n471};
  /* fplog32.vhdl:920:42  */
  assign n473 = n469 == n472;
  /* fplog32.vhdl:920:17  */
  assign n474 = n473 ? 1'b1 : 1'b0;
  /* fplog32.vhdl:921:22  */
  assign n476 = level4_d1[6:0]; // extract
  /* fplog32.vhdl:921:35  */
  assign n477 = digit3_d1 ? n476 : n478;
  /* fplog32.vhdl:921:68  */
  assign n478 = level4_d1[14:8]; // extract
  /* fplog32.vhdl:922:28  */
  assign n480 = level3[6:3]; // extract
  assign n481 = {sozb_d2, sozb_d2, sozb_d2, sozb_d2};
  /* fplog32.vhdl:922:41  */
  assign n482 = n480 == n481;
  /* fplog32.vhdl:922:17  */
  assign n483 = n482 ? 1'b1 : 1'b0;
  /* fplog32.vhdl:923:19  */
  assign n485 = level3[2:0]; // extract
  /* fplog32.vhdl:923:32  */
  assign n486 = digit2 ? n485 : n487;
  /* fplog32.vhdl:923:59  */
  assign n487 = level3[6:4]; // extract
  /* fplog32.vhdl:925:30  */
  assign n488 = ~ozb_d3;
  /* fplog32.vhdl:925:19  */
  assign n489 = n488 ? level2_d1 : n490;
  /* fplog32.vhdl:925:41  */
  assign n490 = ~level2_d1;
  /* fplog32.vhdl:927:12  */
  assign n493 = z == 3'b000;
  /* fplog32.vhdl:928:12  */
  assign n496 = z == 3'b001;
  /* fplog32.vhdl:929:12  */
  assign n499 = z == 3'b010;
  /* fplog32.vhdl:930:12  */
  assign n502 = z == 3'b011;
  assign n504 = {n502, n499, n496, n493};
  /* fplog32.vhdl:926:4  */
  always @*
    case (n504)
      4'b1000: n505 = 2'b01;
      4'b0100: n505 = 2'b01;
      4'b0010: n505 = 2'b10;
      4'b0001: n505 = 2'b11;
      default: n505 = 2'b00;
    endcase
  /* fplog32.vhdl:932:29  */
  assign n506 = {digit4_d2, digit3_d1};
  /* fplog32.vhdl:932:50  */
  assign n507 = {n506, digit2};
  /* fplog32.vhdl:933:24  */
  assign n509 = {outhighbits_d1, lowbits};
  /* fplog32.vhdl:899:10  */
  always @(posedge clk)
    n510 <= sozb;
  /* fplog32.vhdl:899:10  */
  always @(posedge clk)
    n511 <= sozb_d1;
  /* fplog32.vhdl:899:10  */
  always @(posedge clk)
    n512 <= level5;
  /* fplog32.vhdl:899:10  */
  always @(posedge clk)
    n513 <= digit4;
  /* fplog32.vhdl:899:10  */
  always @(posedge clk)
    n514 <= digit4_d1;
  /* fplog32.vhdl:899:10  */
  always @(posedge clk)
    n515 <= level4;
  /* fplog32.vhdl:899:10  */
  always @(posedge clk)
    n516 <= digit3;
  /* fplog32.vhdl:899:10  */
  always @(posedge clk)
    n517 <= level2;
  /* fplog32.vhdl:899:10  */
  always @(posedge clk)
    n518 <= outhighbits;
  /* fplog32.vhdl:899:10  */
  always @(posedge clk)
    n519 <= ozb;
  /* fplog32.vhdl:899:10  */
  always @(posedge clk)
    n520 <= ozb_d1;
  /* fplog32.vhdl:899:10  */
  always @(posedge clk)
    n521 <= ozb_d2;
endmodule

module top_module
  (input  clk,
   input  [33:0] X,
   output [33:0] R);
  wire [2:0] xexnsgn;
  wire [2:0] xexnsgn_d1;
  wire [2:0] xexnsgn_d2;
  wire [2:0] xexnsgn_d3;
  wire [2:0] xexnsgn_d4;
  wire [2:0] xexnsgn_d5;
  wire [2:0] xexnsgn_d6;
  wire [2:0] xexnsgn_d7;
  wire [2:0] xexnsgn_d8;
  wire [2:0] xexnsgn_d9;
  wire [2:0] xexnsgn_d10;
  wire [2:0] xexnsgn_d11;
  wire [2:0] xexnsgn_d12;
  wire firstbit;
  wire [24:0] y0;
  wire [24:0] y0_d1;
  wire [22:0] y0h;
  wire sr;
  wire sr_d1;
  wire sr_d2;
  wire sr_d3;
  wire sr_d4;
  wire sr_d5;
  wire sr_d6;
  wire sr_d7;
  wire sr_d8;
  wire sr_d9;
  wire sr_d10;
  wire sr_d11;
  wire sr_d12;
  wire [11:0] absz0;
  wire [7:0] e;
  wire [7:0] abse;
  wire eeqzero;
  wire eeqzero_d1;
  wire eeqzero_d2;
  wire eeqzero_d3;
  wire eeqzero_d4;
  wire [4:0] lzo;
  wire [4:0] lzo_d1;
  wire [4:0] lzo_d2;
  wire [4:0] lzo_d3;
  wire [4:0] pfinal_s;
  wire [4:0] pfinal_s_d1;
  wire [4:0] pfinal_s_d2;
  wire [4:0] pfinal_s_d3;
  wire [5:0] shiftval;
  wire [3:0] shiftvalinl;
  wire [3:0] shiftvalinr;
  wire dorr;
  wire dorr_d1;
  wire dorr_d2;
  wire \small ;
  wire small_d1;
  wire small_d2;
  wire small_d3;
  wire small_d4;
  wire small_d5;
  wire small_d6;
  wire small_d7;
  wire small_d8;
  wire [23:0] small_absz0_normd_full;
  wire [11:0] small_absz0_normd;
  wire [11:0] small_absz0_normd_d1;
  wire [8:0] a0;
  wire [9:0] inva0;
  wire [9:0] inva0_d1;
  wire [9:0] inva0_copy9;
  wire [34:0] p0;
  wire [25:0] z1;
  wire [6:0] a1;
  wire [6:0] a1_d1;
  wire [18:0] b1;
  wire [25:0] zm1;
  wire [25:0] zm1_d1;
  wire [32:0] p1;
  wire [33:0] y1;
  wire [26:0] eiy1;
  wire [26:0] addxiter1;
  wire [26:0] eiypb1;
  wire [26:0] pp1;
  wire [26:0] z2;
  wire [26:0] zfinal;
  wire [26:0] zfinal_d1;
  wire [26:0] zfinal_d2;
  wire [15:0] squarerin;
  wire [31:0] z2o2_full;
  wire [31:0] z2o2_full_dummy;
  wire [12:0] z2o2_normal;
  wire [26:0] addfinallog1py;
  wire [26:0] log1p_normal;
  wire [39:0] l0;
  wire [39:0] s1;
  wire [32:0] l1;
  wire [32:0] l1_copy23;
  wire [39:0] sopx1;
  wire [39:0] s2;
  wire [39:0] almostlog;
  wire [39:0] adderlogf_normaly;
  wire [39:0] logf_normal;
  wire [34:0] abselog2;
  wire [47:0] abselog2_pad;
  wire [47:0] logf_normal_pad;
  wire [47:0] lnaddx;
  wire [47:0] lnaddy;
  wire [47:0] log_normal;
  wire [39:0] log_normal_normd;
  wire [39:0] log_normal_normd_d1;
  wire [4:0] e_normal;
  wire [15:0] z2o2_small_bs;
  wire [30:0] z2o2_small_s;
  wire [28:0] z2o2_small;
  wire [28:0] z_small;
  wire [28:0] log_smally;
  wire nsrcin;
  wire [28:0] log_small;
  wire [1:0] e0_sub;
  wire ufl;
  wire ufl_d1;
  wire ufl_d2;
  wire ufl_d3;
  wire ufl_d4;
  wire ufl_d5;
  wire ufl_d6;
  wire ufl_d7;
  wire ufl_d8;
  wire ufl_d9;
  wire ufl_d10;
  wire ufl_d11;
  wire ufl_d12;
  wire [7:0] e_small;
  wire [7:0] e_small_d1;
  wire [7:0] e_small_d2;
  wire [7:0] e_small_d3;
  wire [7:0] e_small_d4;
  wire [7:0] e_small_d5;
  wire [26:0] log_small_normd;
  wire [26:0] log_small_normd_d1;
  wire [26:0] log_small_normd_d2;
  wire [26:0] log_small_normd_d3;
  wire [26:0] log_small_normd_d4;
  wire [26:0] log_small_normd_d5;
  wire [26:0] log_small_normd_d6;
  wire [7:0] e0offset;
  wire [7:0] e0offset_d1;
  wire [7:0] e0offset_d2;
  wire [7:0] e0offset_d3;
  wire [7:0] e0offset_d4;
  wire [7:0] e0offset_d5;
  wire [7:0] e0offset_d6;
  wire [7:0] e0offset_d7;
  wire [7:0] e0offset_d8;
  wire [7:0] e0offset_d9;
  wire [7:0] e0offset_d10;
  wire [7:0] e0offset_d11;
  wire [7:0] er;
  wire [26:0] log_g;
  wire round;
  wire [30:0] frax;
  wire [30:0] fray;
  wire [30:0] efr;
  wire [2:0] rexn;
  wire [2:0] n91;
  wire n92;
  wire [22:0] n93;
  wire [23:0] n95;
  wire [24:0] n97;
  wire n98;
  wire [24:0] n99;
  wire [22:0] n100;
  wire [24:0] n102;
  wire [22:0] n103;
  wire [7:0] n105;
  wire n107;
  wire n108;
  wire n109;
  wire n110;
  wire [11:0] n111;
  wire n112;
  wire [11:0] n113;
  wire [11:0] n114;
  wire [11:0] n116;
  wire [7:0] n117;
  wire n118;
  wire [7:0] n120;
  wire [7:0] n121;
  wire [7:0] n123;
  wire [7:0] n124;
  wire n127;
  wire n128;
  wire [4:0] lzoc1_n130;
  wire [5:0] n135;
  wire [5:0] n137;
  wire [5:0] n138;
  wire [3:0] n139;
  wire [3:0] n140;
  wire n141;
  wire n142;
  wire n143;
  wire [23:0] small_lshift_n144;
  wire [11:0] n147;
  wire [8:0] n148;
  wire [9:0] inva0table_n149;
  wire [34:0] n152;
  wire [34:0] n153;
  wire [34:0] n154;
  wire [25:0] n155;
  wire [6:0] n156;
  wire [18:0] n157;
  wire [32:0] n158;
  wire [32:0] n159;
  wire [32:0] n160;
  wire [33:0] n162;
  wire [26:0] n163;
  wire n164;
  wire [26:0] n165;
  wire [25:0] n166;
  wire [26:0] n168;
  wire [19:0] n170;
  wire [26:0] n172;
  localparam n173 = 1'b0;
  wire [26:0] additer1_1_n174;
  wire [25:0] n177;
  wire [25:0] n178;
  wire [26:0] n180;
  localparam n181 = 1'b1;
  wire [26:0] additer2_1_n182;
  wire [15:0] n185;
  wire [15:0] n186;
  wire [15:0] n188;
  wire [31:0] n189;
  wire [31:0] n190;
  wire [31:0] n191;
  wire [12:0] n192;
  wire [12:0] n193;
  wire [26:0] n195;
  localparam n196 = 1'b1;
  wire [26:0] addfinallog1p_normaladder_n197;
  wire [39:0] logtable0_n200;
  wire [32:0] logtable1_n203;
  wire [39:0] n207;
  localparam n208 = 1'b0;
  wire [39:0] adders1_n209;
  wire [39:0] n213;
  localparam n214 = 1'b0;
  wire [39:0] adderlogf_normal_n215;
  wire [34:0] mullog2_n218;
  wire [47:0] n222;
  wire n223;
  wire n224;
  wire n225;
  wire n226;
  wire n227;
  wire n228;
  wire n229;
  wire n230;
  wire [3:0] n231;
  wire [3:0] n232;
  wire [7:0] n233;
  wire [47:0] n234;
  wire n235;
  wire [47:0] n236;
  wire [47:0] n237;
  wire [47:0] lnadder_n238;
  wire [4:0] final_norm_n241;
  wire [39:0] final_norm_n242;
  wire [15:0] n247;
  wire [30:0] ao_rshift_n248;
  wire [15:0] n251;
  wire [28:0] n253;
  wire [28:0] n255;
  wire [28:0] n256;
  wire [28:0] n257;
  wire n258;
  wire [28:0] log_small_adder_n259;
  wire n263;
  wire [1:0] n264;
  wire [1:0] n266;
  wire n268;
  wire [1:0] n269;
  wire [7:0] n273;
  wire [7:0] n275;
  wire [7:0] n276;
  wire [26:0] n277;
  wire n278;
  wire [26:0] n279;
  wire [26:0] n280;
  wire n281;
  wire [26:0] n282;
  wire [26:0] n283;
  wire [7:0] n285;
  wire [7:0] n287;
  wire [7:0] n288;
  wire [25:0] n289;
  wire [26:0] n291;
  wire [26:0] n292;
  wire [26:0] n293;
  wire n294;
  wire [22:0] n295;
  wire [30:0] n296;
  wire [30:0] n298;
  localparam n299 = 1'b0;
  wire [30:0] finalroundadder_n300;
  wire n304;
  wire n305;
  wire n306;
  wire n307;
  wire n308;
  wire n309;
  wire n310;
  wire n311;
  wire n312;
  wire [2:0] n313;
  wire [1:0] n315;
  wire n317;
  wire [2:0] n318;
  wire [1:0] n320;
  wire n322;
  wire [2:0] n323;
  wire [2:0] n325;
  wire n326;
  wire n327;
  wire n328;
  wire n329;
  wire n330;
  wire n331;
  wire n332;
  wire n333;
  wire n334;
  wire n335;
  wire [2:0] n336;
  wire [2:0] n338;
  wire [33:0] n339;
  reg [2:0] n340;
  reg [2:0] n341;
  reg [2:0] n342;
  reg [2:0] n343;
  reg [2:0] n344;
  reg [2:0] n345;
  reg [2:0] n346;
  reg [2:0] n347;
  reg [2:0] n348;
  reg [2:0] n349;
  reg [2:0] n350;
  reg [2:0] n351;
  reg [24:0] n352;
  reg n353;
  reg n354;
  reg n355;
  reg n356;
  reg n357;
  reg n358;
  reg n359;
  reg n360;
  reg n361;
  reg n362;
  reg n363;
  reg n364;
  reg n365;
  reg n366;
  reg n367;
  reg n368;
  reg [4:0] n369;
  reg [4:0] n370;
  reg [4:0] n371;
  reg [4:0] n372;
  reg [4:0] n373;
  reg [4:0] n374;
  reg n375;
  reg n376;
  reg n377;
  reg n378;
  reg n379;
  reg n380;
  reg n381;
  reg n382;
  reg n383;
  reg n384;
  reg [11:0] n385;
  reg [9:0] n386;
  reg [6:0] n387;
  reg [25:0] n388;
  reg [26:0] n389;
  reg [26:0] n390;
  reg [39:0] n391;
  reg n392;
  reg n393;
  reg n394;
  reg n395;
  reg n396;
  reg n397;
  reg n398;
  reg n399;
  reg n400;
  reg n401;
  reg n402;
  reg n403;
  reg [7:0] n404;
  reg [7:0] n405;
  reg [7:0] n406;
  reg [7:0] n407;
  reg [7:0] n408;
  reg [26:0] n409;
  reg [26:0] n410;
  reg [26:0] n411;
  reg [26:0] n412;
  reg [26:0] n413;
  reg [26:0] n414;
  reg [7:0] n415;
  reg [7:0] n416;
  reg [7:0] n417;
  reg [7:0] n418;
  reg [7:0] n419;
  reg [7:0] n420;
  reg [7:0] n421;
  reg [7:0] n422;
  reg [7:0] n423;
  reg [7:0] n424;
  reg [7:0] n425;
  assign R = n339; //(module output)
  /* fplog32.vhdl:2787:8  */
  assign xexnsgn = n91; // (signal)
  /* fplog32.vhdl:2787:17  */
  assign xexnsgn_d1 = n340; // (signal)
  /* fplog32.vhdl:2787:29  */
  assign xexnsgn_d2 = n341; // (signal)
  /* fplog32.vhdl:2787:41  */
  assign xexnsgn_d3 = n342; // (signal)
  /* fplog32.vhdl:2787:53  */
  assign xexnsgn_d4 = n343; // (signal)
  /* fplog32.vhdl:2787:65  */
  assign xexnsgn_d5 = n344; // (signal)
  /* fplog32.vhdl:2787:77  */
  assign xexnsgn_d6 = n345; // (signal)
  /* fplog32.vhdl:2787:89  */
  assign xexnsgn_d7 = n346; // (signal)
  /* fplog32.vhdl:2787:101  */
  assign xexnsgn_d8 = n347; // (signal)
  /* fplog32.vhdl:2787:113  */
  assign xexnsgn_d9 = n348; // (signal)
  /* fplog32.vhdl:2787:125  */
  assign xexnsgn_d10 = n349; // (signal)
  /* fplog32.vhdl:2787:138  */
  assign xexnsgn_d11 = n350; // (signal)
  /* fplog32.vhdl:2787:151  */
  assign xexnsgn_d12 = n351; // (signal)
  /* fplog32.vhdl:2789:8  */
  assign firstbit = n92; // (signal)
  /* fplog32.vhdl:2791:8  */
  assign y0 = n99; // (signal)
  /* fplog32.vhdl:2791:12  */
  assign y0_d1 = n352; // (signal)
  /* fplog32.vhdl:2793:8  */
  assign y0h = n103; // (signal)
  /* fplog32.vhdl:2795:8  */
  assign sr = n108; // (signal)
  /* fplog32.vhdl:2795:12  */
  assign sr_d1 = n353; // (signal)
  /* fplog32.vhdl:2795:19  */
  assign sr_d2 = n354; // (signal)
  /* fplog32.vhdl:2795:26  */
  assign sr_d3 = n355; // (signal)
  /* fplog32.vhdl:2795:33  */
  assign sr_d4 = n356; // (signal)
  /* fplog32.vhdl:2795:40  */
  assign sr_d5 = n357; // (signal)
  /* fplog32.vhdl:2795:47  */
  assign sr_d6 = n358; // (signal)
  /* fplog32.vhdl:2795:54  */
  assign sr_d7 = n359; // (signal)
  /* fplog32.vhdl:2795:61  */
  assign sr_d8 = n360; // (signal)
  /* fplog32.vhdl:2795:68  */
  assign sr_d9 = n361; // (signal)
  /* fplog32.vhdl:2795:75  */
  assign sr_d10 = n362; // (signal)
  /* fplog32.vhdl:2795:83  */
  assign sr_d11 = n363; // (signal)
  /* fplog32.vhdl:2795:91  */
  assign sr_d12 = n364; // (signal)
  /* fplog32.vhdl:2797:8  */
  assign absz0 = n113; // (signal)
  /* fplog32.vhdl:2799:8  */
  assign e = n121; // (signal)
  /* fplog32.vhdl:2801:8  */
  assign abse = n124; // (signal)
  /* fplog32.vhdl:2803:8  */
  assign eeqzero = n128; // (signal)
  /* fplog32.vhdl:2803:17  */
  assign eeqzero_d1 = n365; // (signal)
  /* fplog32.vhdl:2803:29  */
  assign eeqzero_d2 = n366; // (signal)
  /* fplog32.vhdl:2803:41  */
  assign eeqzero_d3 = n367; // (signal)
  /* fplog32.vhdl:2803:53  */
  assign eeqzero_d4 = n368; // (signal)
  /* fplog32.vhdl:2805:8  */
  assign lzo = lzoc1_n130; // (signal)
  /* fplog32.vhdl:2805:13  */
  assign lzo_d1 = n369; // (signal)
  /* fplog32.vhdl:2805:21  */
  assign lzo_d2 = n370; // (signal)
  /* fplog32.vhdl:2805:29  */
  assign lzo_d3 = n371; // (signal)
  /* fplog32.vhdl:2807:8  */
  assign pfinal_s = 5'b01101; // (signal)
  /* fplog32.vhdl:2807:18  */
  assign pfinal_s_d1 = n372; // (signal)
  /* fplog32.vhdl:2807:31  */
  assign pfinal_s_d2 = n373; // (signal)
  /* fplog32.vhdl:2807:44  */
  assign pfinal_s_d3 = n374; // (signal)
  /* fplog32.vhdl:2809:8  */
  assign shiftval = n138; // (signal)
  /* fplog32.vhdl:2811:8  */
  assign shiftvalinl = n139; // (signal)
  /* fplog32.vhdl:2813:8  */
  assign shiftvalinr = n140; // (signal)
  /* fplog32.vhdl:2815:8  */
  assign dorr = n141; // (signal)
  /* fplog32.vhdl:2815:14  */
  assign dorr_d1 = n375; // (signal)
  /* fplog32.vhdl:2815:23  */
  assign dorr_d2 = n376; // (signal)
  /* fplog32.vhdl:2817:8  */
  assign \small  = n143; // (signal)
  /* fplog32.vhdl:2817:15  */
  assign small_d1 = n377; // (signal)
  /* fplog32.vhdl:2817:25  */
  assign small_d2 = n378; // (signal)
  /* fplog32.vhdl:2817:35  */
  assign small_d3 = n379; // (signal)
  /* fplog32.vhdl:2817:45  */
  assign small_d4 = n380; // (signal)
  /* fplog32.vhdl:2817:55  */
  assign small_d5 = n381; // (signal)
  /* fplog32.vhdl:2817:65  */
  assign small_d6 = n382; // (signal)
  /* fplog32.vhdl:2817:75  */
  assign small_d7 = n383; // (signal)
  /* fplog32.vhdl:2817:85  */
  assign small_d8 = n384; // (signal)
  /* fplog32.vhdl:2819:8  */
  assign small_absz0_normd_full = small_lshift_n144; // (signal)
  /* fplog32.vhdl:2821:8  */
  assign small_absz0_normd = n147; // (signal)
  /* fplog32.vhdl:2821:27  */
  assign small_absz0_normd_d1 = n385; // (signal)
  /* fplog32.vhdl:2823:8  */
  assign a0 = n148; // (signal)
  /* fplog32.vhdl:2825:8  */
  assign inva0 = inva0_copy9; // (signal)
  /* fplog32.vhdl:2825:15  */
  assign inva0_d1 = n386; // (signal)
  /* fplog32.vhdl:2827:8  */
  assign inva0_copy9 = inva0table_n149; // (signal)
  /* fplog32.vhdl:2829:8  */
  assign p0 = n154; // (signal)
  /* fplog32.vhdl:2831:8  */
  assign z1 = n155; // (signal)
  /* fplog32.vhdl:2833:8  */
  assign a1 = n156; // (signal)
  /* fplog32.vhdl:2833:12  */
  assign a1_d1 = n387; // (signal)
  /* fplog32.vhdl:2835:8  */
  assign b1 = n157; // (signal)
  /* fplog32.vhdl:2837:8  */
  assign zm1 = z1; // (signal)
  /* fplog32.vhdl:2837:13  */
  assign zm1_d1 = n388; // (signal)
  /* fplog32.vhdl:2839:8  */
  assign p1 = n160; // (signal)
  /* fplog32.vhdl:2841:8  */
  assign y1 = n162; // (signal)
  /* fplog32.vhdl:2843:8  */
  assign eiy1 = n165; // (signal)
  /* fplog32.vhdl:2845:8  */
  assign addxiter1 = n172; // (signal)
  /* fplog32.vhdl:2847:8  */
  assign eiypb1 = additer1_1_n174; // (signal)
  /* fplog32.vhdl:2849:8  */
  assign pp1 = n180; // (signal)
  /* fplog32.vhdl:2851:8  */
  assign z2 = additer2_1_n182; // (signal)
  /* fplog32.vhdl:2853:8  */
  assign zfinal = z2; // (signal)
  /* fplog32.vhdl:2853:16  */
  assign zfinal_d1 = n389; // (signal)
  /* fplog32.vhdl:2853:27  */
  assign zfinal_d2 = n390; // (signal)
  /* fplog32.vhdl:2855:8  */
  assign squarerin = n186; // (signal)
  /* fplog32.vhdl:2857:8  */
  assign z2o2_full = n191; // (signal)
  /* fplog32.vhdl:2859:8  */
  assign z2o2_full_dummy = z2o2_full; // (signal)
  /* fplog32.vhdl:2861:8  */
  assign z2o2_normal = n192; // (signal)
  /* fplog32.vhdl:2863:8  */
  assign addfinallog1py = n195; // (signal)
  /* fplog32.vhdl:2865:8  */
  assign log1p_normal = addfinallog1p_normaladder_n197; // (signal)
  /* fplog32.vhdl:2867:8  */
  assign l0 = logtable0_n200; // (signal)
  /* fplog32.vhdl:2869:8  */
  assign s1 = l0; // (signal)
  /* fplog32.vhdl:2871:8  */
  assign l1 = l1_copy23; // (signal)
  /* fplog32.vhdl:2873:8  */
  assign l1_copy23 = logtable1_n203; // (signal)
  /* fplog32.vhdl:2875:8  */
  assign sopx1 = n207; // (signal)
  /* fplog32.vhdl:2877:8  */
  assign s2 = adders1_n209; // (signal)
  /* fplog32.vhdl:2879:8  */
  assign almostlog = s2; // (signal)
  /* fplog32.vhdl:2881:8  */
  assign adderlogf_normaly = n213; // (signal)
  /* fplog32.vhdl:2883:8  */
  assign logf_normal = adderlogf_normal_n215; // (signal)
  /* fplog32.vhdl:2885:8  */
  assign abselog2 = mullog2_n218; // (signal)
  /* fplog32.vhdl:2887:8  */
  assign abselog2_pad = n222; // (signal)
  /* fplog32.vhdl:2889:8  */
  assign logf_normal_pad = n234; // (signal)
  /* fplog32.vhdl:2891:8  */
  assign lnaddx = abselog2_pad; // (signal)
  /* fplog32.vhdl:2893:8  */
  assign lnaddy = n236; // (signal)
  /* fplog32.vhdl:2895:8  */
  assign log_normal = lnadder_n238; // (signal)
  /* fplog32.vhdl:2897:8  */
  assign log_normal_normd = final_norm_n242; // (signal)
  /* fplog32.vhdl:2897:26  */
  assign log_normal_normd_d1 = n391; // (signal)
  /* fplog32.vhdl:2899:8  */
  assign e_normal = final_norm_n241; // (signal)
  /* fplog32.vhdl:2901:8  */
  assign z2o2_small_bs = n247; // (signal)
  /* fplog32.vhdl:2903:8  */
  assign z2o2_small_s = ao_rshift_n248; // (signal)
  /* fplog32.vhdl:2905:8  */
  assign z2o2_small = n253; // (signal)
  /* fplog32.vhdl:2907:8  */
  assign z_small = n255; // (signal)
  /* fplog32.vhdl:2909:8  */
  assign log_smally = n256; // (signal)
  /* fplog32.vhdl:2911:8  */
  assign nsrcin = n258; // (signal)
  /* fplog32.vhdl:2913:8  */
  assign log_small = log_small_adder_n259; // (signal)
  /* fplog32.vhdl:2915:8  */
  assign e0_sub = n264; // (signal)
  /* fplog32.vhdl:2917:8  */
  assign ufl = 1'b0; // (signal)
  /* fplog32.vhdl:2917:13  */
  assign ufl_d1 = n392; // (signal)
  /* fplog32.vhdl:2917:21  */
  assign ufl_d2 = n393; // (signal)
  /* fplog32.vhdl:2917:29  */
  assign ufl_d3 = n394; // (signal)
  /* fplog32.vhdl:2917:37  */
  assign ufl_d4 = n395; // (signal)
  /* fplog32.vhdl:2917:45  */
  assign ufl_d5 = n396; // (signal)
  /* fplog32.vhdl:2917:53  */
  assign ufl_d6 = n397; // (signal)
  /* fplog32.vhdl:2917:61  */
  assign ufl_d7 = n398; // (signal)
  /* fplog32.vhdl:2917:69  */
  assign ufl_d8 = n399; // (signal)
  /* fplog32.vhdl:2917:77  */
  assign ufl_d9 = n400; // (signal)
  /* fplog32.vhdl:2917:85  */
  assign ufl_d10 = n401; // (signal)
  /* fplog32.vhdl:2917:94  */
  assign ufl_d11 = n402; // (signal)
  /* fplog32.vhdl:2917:103  */
  assign ufl_d12 = n403; // (signal)
  /* fplog32.vhdl:2919:8  */
  assign e_small = n276; // (signal)
  /* fplog32.vhdl:2919:17  */
  assign e_small_d1 = n404; // (signal)
  /* fplog32.vhdl:2919:29  */
  assign e_small_d2 = n405; // (signal)
  /* fplog32.vhdl:2919:41  */
  assign e_small_d3 = n406; // (signal)
  /* fplog32.vhdl:2919:53  */
  assign e_small_d4 = n407; // (signal)
  /* fplog32.vhdl:2919:65  */
  assign e_small_d5 = n408; // (signal)
  /* fplog32.vhdl:2921:8  */
  assign log_small_normd = n279; // (signal)
  /* fplog32.vhdl:2921:25  */
  assign log_small_normd_d1 = n409; // (signal)
  /* fplog32.vhdl:2921:45  */
  assign log_small_normd_d2 = n410; // (signal)
  /* fplog32.vhdl:2921:65  */
  assign log_small_normd_d3 = n411; // (signal)
  /* fplog32.vhdl:2921:85  */
  assign log_small_normd_d4 = n412; // (signal)
  /* fplog32.vhdl:2921:105  */
  assign log_small_normd_d5 = n413; // (signal)
  /* fplog32.vhdl:2921:125  */
  assign log_small_normd_d6 = n414; // (signal)
  /* fplog32.vhdl:2923:8  */
  assign e0offset = 8'b10000110; // (signal)
  /* fplog32.vhdl:2923:18  */
  assign e0offset_d1 = n415; // (signal)
  /* fplog32.vhdl:2923:31  */
  assign e0offset_d2 = n416; // (signal)
  /* fplog32.vhdl:2923:44  */
  assign e0offset_d3 = n417; // (signal)
  /* fplog32.vhdl:2923:57  */
  assign e0offset_d4 = n418; // (signal)
  /* fplog32.vhdl:2923:70  */
  assign e0offset_d5 = n419; // (signal)
  /* fplog32.vhdl:2923:83  */
  assign e0offset_d6 = n420; // (signal)
  /* fplog32.vhdl:2923:96  */
  assign e0offset_d7 = n421; // (signal)
  /* fplog32.vhdl:2923:109  */
  assign e0offset_d8 = n422; // (signal)
  /* fplog32.vhdl:2923:122  */
  assign e0offset_d9 = n423; // (signal)
  /* fplog32.vhdl:2923:135  */
  assign e0offset_d10 = n424; // (signal)
  /* fplog32.vhdl:2923:149  */
  assign e0offset_d11 = n425; // (signal)
  /* fplog32.vhdl:2925:8  */
  assign er = n285; // (signal)
  /* fplog32.vhdl:2927:8  */
  assign log_g = n292; // (signal)
  /* fplog32.vhdl:2929:8  */
  assign round = n294; // (signal)
  /* fplog32.vhdl:2931:8  */
  assign frax = n296; // (signal)
  /* fplog32.vhdl:2933:8  */
  assign fray = n298; // (signal)
  /* fplog32.vhdl:2935:8  */
  assign efr = finalroundadder_n300; // (signal)
  /* fplog32.vhdl:2937:8  */
  assign rexn = n313; // (signal)
  /* fplog32.vhdl:3038:17  */
  assign n91 = X[33:31]; // extract
  /* fplog32.vhdl:3039:18  */
  assign n92 = X[22]; // extract
  /* fplog32.vhdl:3040:17  */
  assign n93 = X[22:0]; // extract
  /* fplog32.vhdl:3040:14  */
  assign n95 = {1'b1, n93};
  /* fplog32.vhdl:3040:33  */
  assign n97 = {n95, 1'b0};
  /* fplog32.vhdl:3040:53  */
  assign n98 = ~firstbit;
  /* fplog32.vhdl:3040:39  */
  assign n99 = n98 ? n97 : n102;
  /* fplog32.vhdl:3040:72  */
  assign n100 = X[22:0]; // extract
  /* fplog32.vhdl:3040:69  */
  assign n102 = {2'b01, n100};
  /* fplog32.vhdl:3041:13  */
  assign n103 = y0[23:1]; // extract
  /* fplog32.vhdl:3043:24  */
  assign n105 = X[30:23]; // extract
  /* fplog32.vhdl:3043:44  */
  assign n107 = n105 == 8'b01111111;
  /* fplog32.vhdl:3043:16  */
  assign n108 = n107 ? 1'b0 : n110;
  /* fplog32.vhdl:3044:16  */
  assign n109 = X[30]; // extract
  /* fplog32.vhdl:3044:11  */
  assign n110 = ~n109;
  /* fplog32.vhdl:3045:17  */
  assign n111 = y0[11:0]; // extract
  /* fplog32.vhdl:3045:57  */
  assign n112 = ~sr;
  /* fplog32.vhdl:3045:49  */
  assign n113 = n112 ? n111 : n116;
  /* fplog32.vhdl:3046:49  */
  assign n114 = y0[11:0]; // extract
  /* fplog32.vhdl:3046:45  */
  assign n116 = 12'b000000000000 - n114;
  /* fplog32.vhdl:3047:11  */
  assign n117 = X[30:23]; // extract
  /* fplog32.vhdl:3047:67  */
  assign n118 = ~firstbit;
  /* fplog32.vhdl:3047:64  */
  assign n120 = {7'b0111111, n118};
  /* fplog32.vhdl:3047:32  */
  assign n121 = n117 - n120;
  /* fplog32.vhdl:3048:36  */
  assign n123 = 8'b00000000 - e;
  /* fplog32.vhdl:3048:43  */
  assign n124 = sr ? n123 : e;
  /* fplog32.vhdl:3049:25  */
  assign n127 = e == 8'b00000000;
  /* fplog32.vhdl:3049:19  */
  assign n128 = n127 ? 1'b1 : 1'b0;
  /* fplog32.vhdl:3050:4  */
  lzoc_23_freq500_uid4 lzoc1 (
    .clk(clk),
    .i(y0h),
    .ozb(firstbit),
    .o(lzoc1_n130));
  /* fplog32.vhdl:3056:21  */
  assign n135 = {1'b0, lzo};
  /* fplog32.vhdl:3056:35  */
  assign n137 = {1'b0, pfinal_s_d3};
  /* fplog32.vhdl:3056:28  */
  assign n138 = n135 - n137;
  /* fplog32.vhdl:3057:27  */
  assign n139 = shiftval[3:0]; // extract
  /* fplog32.vhdl:3058:27  */
  assign n140 = shiftval[3:0]; // extract
  /* fplog32.vhdl:3059:20  */
  assign n141 = shiftval[5]; // extract
  /* fplog32.vhdl:3060:28  */
  assign n142 = ~dorr_d1;
  /* fplog32.vhdl:3060:24  */
  assign n143 = eeqzero_d4 & n142;
  /* fplog32.vhdl:3062:4  */
  leftshifter12_by_max_12_freq500_uid6 small_lshift (
    .clk(clk),
    .x(absz0),
    .s(shiftvalinl),
    .r(small_lshift_n144));
  /* fplog32.vhdl:3067:47  */
  assign n147 = small_absz0_normd_full[11:0]; // extract
  /* fplog32.vhdl:3069:11  */
  assign n148 = X[22:14]; // extract
  /* fplog32.vhdl:3071:4  */
  inva0table_freq500_uid8 inva0table (
    .x(a0),
    .y(inva0table_n149));
  /* fplog32.vhdl:3075:19  */
  assign n152 = {25'b0, inva0_d1};  //  uext
  /* fplog32.vhdl:3075:19  */
  assign n153 = {10'b0, y0_d1};  //  uext
  /* fplog32.vhdl:3075:19  */
  assign n154 = n152 * n153; // umul
  /* fplog32.vhdl:3077:12  */
  assign n155 = p0[25:0]; // extract
  /* fplog32.vhdl:3079:12  */
  assign n156 = z1[25:19]; // extract
  /* fplog32.vhdl:3080:12  */
  assign n157 = z1[18:0]; // extract
  /* fplog32.vhdl:3082:15  */
  assign n158 = {26'b0, a1_d1};  //  uext
  /* fplog32.vhdl:3082:15  */
  assign n159 = {7'b0, zm1_d1};  //  uext
  /* fplog32.vhdl:3082:15  */
  assign n160 = n158 * n159; // umul
  /* fplog32.vhdl:3083:36  */
  assign n162 = {8'b10000000, z1};
  /* fplog32.vhdl:3084:14  */
  assign n163 = y1[33:7]; // extract
  /* fplog32.vhdl:3084:36  */
  assign n164 = a1[6]; // extract
  /* fplog32.vhdl:3084:29  */
  assign n165 = n164 ? n163 : n168;
  /* fplog32.vhdl:3085:20  */
  assign n166 = y1[33:8]; // extract
  /* fplog32.vhdl:3085:16  */
  assign n168 = {1'b0, n166};
  /* fplog32.vhdl:3086:21  */
  assign n170 = {1'b0, b1};
  /* fplog32.vhdl:3086:26  */
  assign n172 = {n170, 7'b0000000};
  /* fplog32.vhdl:3087:4  */
  intadder_27_freq500_uid12 additer1_1 (
    .clk(clk),
    .x(addxiter1),
    .y(eiy1),
    .cin(n173),
    .r(additer1_1_n174));
  /* fplog32.vhdl:3093:39  */
  assign n177 = p1[32:7]; // extract
  /* fplog32.vhdl:3093:33  */
  assign n178 = ~n177;
  /* fplog32.vhdl:3093:31  */
  assign n180 = {1'b1, n178};
  /* fplog32.vhdl:3094:4  */
  intadder_27_freq500_uid15 additer2_1 (
    .clk(clk),
    .x(eiypb1),
    .y(pp1),
    .cin(n181),
    .r(additer2_1_n182));
  /* fplog32.vhdl:3101:26  */
  assign n185 = zfinal_d2[26:11]; // extract
  /* fplog32.vhdl:3101:54  */
  assign n186 = dorr_d2 ? n185 : n188;
  /* fplog32.vhdl:3102:48  */
  assign n188 = {small_absz0_normd_d1, 4'b0000};
  /* fplog32.vhdl:3103:26  */
  assign n189 = {16'b0, squarerin};  //  uext
  /* fplog32.vhdl:3103:26  */
  assign n190 = {16'b0, squarerin};  //  uext
  /* fplog32.vhdl:3103:26  */
  assign n191 = n189 * n190; // umul
  /* fplog32.vhdl:3105:35  */
  assign n192 = z2o2_full_dummy[31:19]; // extract
  /* fplog32.vhdl:3106:50  */
  assign n193 = ~z2o2_normal;
  /* fplog32.vhdl:3106:48  */
  assign n195 = {14'b11111111111111, n193};
  /* fplog32.vhdl:3107:4  */
  intadder_27_freq500_uid18 addfinallog1p_normaladder (
    .clk(clk),
    .x(zfinal),
    .y(addfinallog1py),
    .cin(n196),
    .r(addfinallog1p_normaladder_n197));
  /* fplog32.vhdl:3115:4  */
  logtable0_freq500_uid20 logtable0 (
    .clk(clk),
    .x(a0),
    .y(logtable0_n200));
  /* fplog32.vhdl:3120:4  */
  logtable1_freq500_uid22 logtable1 (
    .x(a1),
    .y(logtable1_n203));
  /* fplog32.vhdl:3124:36  */
  assign n207 = {7'b0000000, l1};
  /* fplog32.vhdl:3125:4  */
  intadder_40_freq500_uid26 adders1 (
    .clk(clk),
    .x(s1),
    .y(sopx1),
    .cin(n208),
    .r(adders1_n209));
  /* fplog32.vhdl:3132:62  */
  assign n213 = {13'b0000000000000, log1p_normal};
  /* fplog32.vhdl:3133:4  */
  intadder_40_freq500_uid29 adderlogf_normal (
    .clk(clk),
    .x(almostlog),
    .y(adderlogf_normaly),
    .cin(n214),
    .r(adderlogf_normal_n215));
  /* fplog32.vhdl:3139:4  */
  fixrealkcm_freq500_uid31 mullog2 (
    .clk(clk),
    .x(abse),
    .r(mullog2_n218));
  /* fplog32.vhdl:3143:31  */
  assign n222 = {abselog2, 13'b0000000000000};
  /* fplog32.vhdl:3144:53  */
  assign n223 = logf_normal[39]; // extract
  /* fplog32.vhdl:3144:53  */
  assign n224 = logf_normal[39]; // extract
  /* fplog32.vhdl:3144:53  */
  assign n225 = logf_normal[39]; // extract
  /* fplog32.vhdl:3144:53  */
  assign n226 = logf_normal[39]; // extract
  /* fplog32.vhdl:3144:53  */
  assign n227 = logf_normal[39]; // extract
  /* fplog32.vhdl:3144:53  */
  assign n228 = logf_normal[39]; // extract
  /* fplog32.vhdl:3144:53  */
  assign n229 = logf_normal[39]; // extract
  /* fplog32.vhdl:3144:53  */
  assign n230 = logf_normal[39]; // extract
  assign n231 = {n230, n229, n228, n227};
  assign n232 = {n226, n225, n224, n223};
  assign n233 = {n231, n232};
  /* fplog32.vhdl:3144:70  */
  assign n234 = {n233, logf_normal};
  /* fplog32.vhdl:3146:40  */
  assign n235 = ~sr_d7;
  /* fplog32.vhdl:3146:30  */
  assign n236 = n235 ? logf_normal_pad : n237;
  /* fplog32.vhdl:3146:50  */
  assign n237 = ~logf_normal_pad;
  /* fplog32.vhdl:3147:4  */
  intadder_48_freq500_uid43 lnadder (
    .clk(clk),
    .x(lnaddx),
    .y(lnaddy),
    .cin(sr),
    .r(lnadder_n238));
  /* fplog32.vhdl:3153:4  */
  normalizer_z_48_40_19_freq500_uid45 final_norm (
    .clk(clk),
    .x(log_normal),
    .count(final_norm_n241),
    .r(final_norm_n242));
  /* fplog32.vhdl:3158:36  */
  assign n247 = z2o2_full_dummy[31:16]; // extract
  /* fplog32.vhdl:3159:4  */
  rightshifter16_by_max_15_freq500_uid47 ao_rshift (
    .clk(clk),
    .x(z2o2_small_bs),
    .s(shiftvalinr),
    .r(ao_rshift_n248));
  /* fplog32.vhdl:3165:61  */
  assign n251 = z2o2_small_s[30:15]; // extract
  /* fplog32.vhdl:3165:47  */
  assign n253 = {13'b0000000000000, n251};
  /* fplog32.vhdl:3167:33  */
  assign n255 = {small_absz0_normd, 17'b00000000000000000};
  /* fplog32.vhdl:3168:29  */
  assign n256 = sr_d6 ? z2o2_small : n257;
  /* fplog32.vhdl:3168:49  */
  assign n257 = ~z2o2_small;
  /* fplog32.vhdl:3169:14  */
  assign n258 = ~sr;
  /* fplog32.vhdl:3170:4  */
  intadder_29_freq500_uid49 log_small_adder (
    .clk(clk),
    .x(z_small),
    .y(log_smally),
    .cin(nsrcin),
    .r(log_small_adder_n259));
  /* fplog32.vhdl:3177:35  */
  assign n263 = log_small[28]; // extract
  /* fplog32.vhdl:3177:21  */
  assign n264 = n263 ? 2'b11 : n269;
  /* fplog32.vhdl:3178:35  */
  assign n266 = log_small[28:27]; // extract
  /* fplog32.vhdl:3178:56  */
  assign n268 = n266 == 2'b01;
  /* fplog32.vhdl:3178:11  */
  assign n269 = n268 ? 2'b10 : 2'b01;
  /* fplog32.vhdl:3184:46  */
  assign n273 = {6'b011111, e0_sub};
  /* fplog32.vhdl:3184:84  */
  assign n275 = {3'b000, lzo_d3};
  /* fplog32.vhdl:3184:57  */
  assign n276 = n273 - n275;
  /* fplog32.vhdl:3185:32  */
  assign n277 = log_small[28:2]; // extract
  /* fplog32.vhdl:3185:64  */
  assign n278 = log_small[28]; // extract
  /* fplog32.vhdl:3185:50  */
  assign n279 = n278 ? n277 : n282;
  /* fplog32.vhdl:3186:26  */
  assign n280 = log_small[27:1]; // extract
  /* fplog32.vhdl:3186:57  */
  assign n281 = log_small[27]; // extract
  /* fplog32.vhdl:3186:12  */
  assign n282 = n281 ? n280 : n283;
  /* fplog32.vhdl:3187:26  */
  assign n283 = log_small[26:0]; // extract
  /* fplog32.vhdl:3189:33  */
  assign n285 = small_d7 ? e_small_d5 : n288;
  /* fplog32.vhdl:3190:48  */
  assign n287 = {3'b000, e_normal};
  /* fplog32.vhdl:3190:25  */
  assign n288 = e0offset_d11 - n287;
  /* fplog32.vhdl:3191:32  */
  assign n289 = log_small_normd_d5[25:0]; // extract
  /* fplog32.vhdl:3191:50  */
  assign n291 = {n289, 1'b0};
  /* fplog32.vhdl:3191:56  */
  assign n292 = small_d7 ? n291 : n293;
  /* fplog32.vhdl:3192:28  */
  assign n293 = log_normal_normd[38:12]; // extract
  /* fplog32.vhdl:3193:18  */
  assign n294 = log_g[3]; // extract
  /* fplog32.vhdl:3195:23  */
  assign n295 = log_g[26:4]; // extract
  /* fplog32.vhdl:3195:16  */
  assign n296 = {er, n295};
  /* fplog32.vhdl:3196:39  */
  assign n298 = {30'b000000000000000000000000000000, round};
  /* fplog32.vhdl:3197:4  */
  intadder_31_freq500_uid52 finalroundadder (
    .clk(clk),
    .x(frax),
    .y(fray),
    .cin(n299),
    .r(finalroundadder_n300));
  /* fplog32.vhdl:3203:36  */
  assign n304 = xexnsgn_d12[2]; // extract
  /* fplog32.vhdl:3203:56  */
  assign n305 = xexnsgn_d12[1]; // extract
  /* fplog32.vhdl:3203:74  */
  assign n306 = xexnsgn_d12[0]; // extract
  /* fplog32.vhdl:3203:60  */
  assign n307 = n305 | n306;
  /* fplog32.vhdl:3203:40  */
  assign n308 = n304 & n307;
  /* fplog32.vhdl:3203:95  */
  assign n309 = xexnsgn_d12[1]; // extract
  /* fplog32.vhdl:3203:114  */
  assign n310 = xexnsgn_d12[0]; // extract
  /* fplog32.vhdl:3203:99  */
  assign n311 = n309 & n310;
  /* fplog32.vhdl:3203:80  */
  assign n312 = n308 | n311;
  /* fplog32.vhdl:3203:18  */
  assign n313 = n312 ? 3'b110 : n318;
  /* fplog32.vhdl:3204:53  */
  assign n315 = xexnsgn_d12[2:1]; // extract
  /* fplog32.vhdl:3204:66  */
  assign n317 = n315 == 2'b00;
  /* fplog32.vhdl:3203:126  */
  assign n318 = n317 ? 3'b101 : n323;
  /* fplog32.vhdl:3205:53  */
  assign n320 = xexnsgn_d12[2:1]; // extract
  /* fplog32.vhdl:3205:66  */
  assign n322 = n320 == 2'b10;
  /* fplog32.vhdl:3204:74  */
  assign n323 = n322 ? 3'b100 : n336;
  /* fplog32.vhdl:3206:36  */
  assign n325 = {2'b00, sr_d12};
  /* fplog32.vhdl:3206:72  */
  assign n326 = log_normal_normd_d1[39]; // extract
  /* fplog32.vhdl:3206:86  */
  assign n327 = ~n326;
  /* fplog32.vhdl:3206:105  */
  assign n328 = ~small_d8;
  /* fplog32.vhdl:3206:92  */
  assign n329 = n328 & n327;
  /* fplog32.vhdl:3206:137  */
  assign n330 = log_small_normd_d6[26]; // extract
  /* fplog32.vhdl:3206:145  */
  assign n331 = ~n330;
  /* fplog32.vhdl:3206:151  */
  assign n332 = small_d8 & n331;
  /* fplog32.vhdl:3206:112  */
  assign n333 = n329 | n332;
  /* fplog32.vhdl:3206:190  */
  assign n334 = small_d8 & ufl_d12;
  /* fplog32.vhdl:3206:172  */
  assign n335 = n333 | n334;
  /* fplog32.vhdl:3205:74  */
  assign n336 = n335 ? n325 : n338;
  /* fplog32.vhdl:3207:37  */
  assign n338 = {2'b01, sr_d12};
  /* fplog32.vhdl:3208:14  */
  assign n339 = {rexn, efr};
  /* fplog32.vhdl:2949:10  */
  always @(posedge clk)
    n340 <= xexnsgn;
  /* fplog32.vhdl:2949:10  */
  always @(posedge clk)
    n341 <= xexnsgn_d1;
  /* fplog32.vhdl:2949:10  */
  always @(posedge clk)
    n342 <= xexnsgn_d2;
  /* fplog32.vhdl:2949:10  */
  always @(posedge clk)
    n343 <= xexnsgn_d3;
  /* fplog32.vhdl:2949:10  */
  always @(posedge clk)
    n344 <= xexnsgn_d4;
  /* fplog32.vhdl:2949:10  */
  always @(posedge clk)
    n345 <= xexnsgn_d5;
  /* fplog32.vhdl:2949:10  */
  always @(posedge clk)
    n346 <= xexnsgn_d6;
  /* fplog32.vhdl:2949:10  */
  always @(posedge clk)
    n347 <= xexnsgn_d7;
  /* fplog32.vhdl:2949:10  */
  always @(posedge clk)
    n348 <= xexnsgn_d8;
  /* fplog32.vhdl:2949:10  */
  always @(posedge clk)
    n349 <= xexnsgn_d9;
  /* fplog32.vhdl:2949:10  */
  always @(posedge clk)
    n350 <= xexnsgn_d10;
  /* fplog32.vhdl:2949:10  */
  always @(posedge clk)
    n351 <= xexnsgn_d11;
  /* fplog32.vhdl:2949:10  */
  always @(posedge clk)
    n352 <= y0;
  /* fplog32.vhdl:2949:10  */
  always @(posedge clk)
    n353 <= sr;
  /* fplog32.vhdl:2949:10  */
  always @(posedge clk)
    n354 <= sr_d1;
  /* fplog32.vhdl:2949:10  */
  always @(posedge clk)
    n355 <= sr_d2;
  /* fplog32.vhdl:2949:10  */
  always @(posedge clk)
    n356 <= sr_d3;
  /* fplog32.vhdl:2949:10  */
  always @(posedge clk)
    n357 <= sr_d4;
  /* fplog32.vhdl:2949:10  */
  always @(posedge clk)
    n358 <= sr_d5;
  /* fplog32.vhdl:2949:10  */
  always @(posedge clk)
    n359 <= sr_d6;
  /* fplog32.vhdl:2949:10  */
  always @(posedge clk)
    n360 <= sr_d7;
  /* fplog32.vhdl:2949:10  */
  always @(posedge clk)
    n361 <= sr_d8;
  /* fplog32.vhdl:2949:10  */
  always @(posedge clk)
    n362 <= sr_d9;
  /* fplog32.vhdl:2949:10  */
  always @(posedge clk)
    n363 <= sr_d10;
  /* fplog32.vhdl:2949:10  */
  always @(posedge clk)
    n364 <= sr_d11;
  /* fplog32.vhdl:2949:10  */
  always @(posedge clk)
    n365 <= eeqzero;
  /* fplog32.vhdl:2949:10  */
  always @(posedge clk)
    n366 <= eeqzero_d1;
  /* fplog32.vhdl:2949:10  */
  always @(posedge clk)
    n367 <= eeqzero_d2;
  /* fplog32.vhdl:2949:10  */
  always @(posedge clk)
    n368 <= eeqzero_d3;
  /* fplog32.vhdl:2949:10  */
  always @(posedge clk)
    n369 <= lzo;
  /* fplog32.vhdl:2949:10  */
  always @(posedge clk)
    n370 <= lzo_d1;
  /* fplog32.vhdl:2949:10  */
  always @(posedge clk)
    n371 <= lzo_d2;
  /* fplog32.vhdl:2949:10  */
  always @(posedge clk)
    n372 <= pfinal_s;
  /* fplog32.vhdl:2949:10  */
  always @(posedge clk)
    n373 <= pfinal_s_d1;
  /* fplog32.vhdl:2949:10  */
  always @(posedge clk)
    n374 <= pfinal_s_d2;
  /* fplog32.vhdl:2949:10  */
  always @(posedge clk)
    n375 <= dorr;
  /* fplog32.vhdl:2949:10  */
  always @(posedge clk)
    n376 <= dorr_d1;
  /* fplog32.vhdl:2949:10  */
  always @(posedge clk)
    n377 <= \small ;
  /* fplog32.vhdl:2949:10  */
  always @(posedge clk)
    n378 <= small_d1;
  /* fplog32.vhdl:2949:10  */
  always @(posedge clk)
    n379 <= small_d2;
  /* fplog32.vhdl:2949:10  */
  always @(posedge clk)
    n380 <= small_d3;
  /* fplog32.vhdl:2949:10  */
  always @(posedge clk)
    n381 <= small_d4;
  /* fplog32.vhdl:2949:10  */
  always @(posedge clk)
    n382 <= small_d5;
  /* fplog32.vhdl:2949:10  */
  always @(posedge clk)
    n383 <= small_d6;
  /* fplog32.vhdl:2949:10  */
  always @(posedge clk)
    n384 <= small_d7;
  /* fplog32.vhdl:2949:10  */
  always @(posedge clk)
    n385 <= small_absz0_normd;
  /* fplog32.vhdl:2949:10  */
  always @(posedge clk)
    n386 <= inva0;
  /* fplog32.vhdl:2949:10  */
  always @(posedge clk)
    n387 <= a1;
  /* fplog32.vhdl:2949:10  */
  always @(posedge clk)
    n388 <= zm1;
  /* fplog32.vhdl:2949:10  */
  always @(posedge clk)
    n389 <= zfinal;
  /* fplog32.vhdl:2949:10  */
  always @(posedge clk)
    n390 <= zfinal_d1;
  /* fplog32.vhdl:2949:10  */
  always @(posedge clk)
    n391 <= log_normal_normd;
  /* fplog32.vhdl:2949:10  */
  always @(posedge clk)
    n392 <= ufl;
  /* fplog32.vhdl:2949:10  */
  always @(posedge clk)
    n393 <= ufl_d1;
  /* fplog32.vhdl:2949:10  */
  always @(posedge clk)
    n394 <= ufl_d2;
  /* fplog32.vhdl:2949:10  */
  always @(posedge clk)
    n395 <= ufl_d3;
  /* fplog32.vhdl:2949:10  */
  always @(posedge clk)
    n396 <= ufl_d4;
  /* fplog32.vhdl:2949:10  */
  always @(posedge clk)
    n397 <= ufl_d5;
  /* fplog32.vhdl:2949:10  */
  always @(posedge clk)
    n398 <= ufl_d6;
  /* fplog32.vhdl:2949:10  */
  always @(posedge clk)
    n399 <= ufl_d7;
  /* fplog32.vhdl:2949:10  */
  always @(posedge clk)
    n400 <= ufl_d8;
  /* fplog32.vhdl:2949:10  */
  always @(posedge clk)
    n401 <= ufl_d9;
  /* fplog32.vhdl:2949:10  */
  always @(posedge clk)
    n402 <= ufl_d10;
  /* fplog32.vhdl:2949:10  */
  always @(posedge clk)
    n403 <= ufl_d11;
  /* fplog32.vhdl:2949:10  */
  always @(posedge clk)
    n404 <= e_small;
  /* fplog32.vhdl:2949:10  */
  always @(posedge clk)
    n405 <= e_small_d1;
  /* fplog32.vhdl:2949:10  */
  always @(posedge clk)
    n406 <= e_small_d2;
  /* fplog32.vhdl:2949:10  */
  always @(posedge clk)
    n407 <= e_small_d3;
  /* fplog32.vhdl:2949:10  */
  always @(posedge clk)
    n408 <= e_small_d4;
  /* fplog32.vhdl:2949:10  */
  always @(posedge clk)
    n409 <= log_small_normd;
  /* fplog32.vhdl:2949:10  */
  always @(posedge clk)
    n410 <= log_small_normd_d1;
  /* fplog32.vhdl:2949:10  */
  always @(posedge clk)
    n411 <= log_small_normd_d2;
  /* fplog32.vhdl:2949:10  */
  always @(posedge clk)
    n412 <= log_small_normd_d3;
  /* fplog32.vhdl:2949:10  */
  always @(posedge clk)
    n413 <= log_small_normd_d4;
  /* fplog32.vhdl:2949:10  */
  always @(posedge clk)
    n414 <= log_small_normd_d5;
  /* fplog32.vhdl:2949:10  */
  always @(posedge clk)
    n415 <= e0offset;
  /* fplog32.vhdl:2949:10  */
  always @(posedge clk)
    n416 <= e0offset_d1;
  /* fplog32.vhdl:2949:10  */
  always @(posedge clk)
    n417 <= e0offset_d2;
  /* fplog32.vhdl:2949:10  */
  always @(posedge clk)
    n418 <= e0offset_d3;
  /* fplog32.vhdl:2949:10  */
  always @(posedge clk)
    n419 <= e0offset_d4;
  /* fplog32.vhdl:2949:10  */
  always @(posedge clk)
    n420 <= e0offset_d5;
  /* fplog32.vhdl:2949:10  */
  always @(posedge clk)
    n421 <= e0offset_d6;
  /* fplog32.vhdl:2949:10  */
  always @(posedge clk)
    n422 <= e0offset_d7;
  /* fplog32.vhdl:2949:10  */
  always @(posedge clk)
    n423 <= e0offset_d8;
  /* fplog32.vhdl:2949:10  */
  always @(posedge clk)
    n424 <= e0offset_d9;
  /* fplog32.vhdl:2949:10  */
  always @(posedge clk)
    n425 <= e0offset_d10;
endmodule

