module fixrealkcm_freq500_uid84_t0_freq500_uid87
  (input  [4:0] x,
   output [17:0] y);
  wire [17:0] y0;
  wire [17:0] y1;
  wire n6559;
  wire n6562;
  wire n6565;
  wire n6568;
  wire n6571;
  wire n6574;
  wire n6577;
  wire n6580;
  wire n6583;
  wire n6586;
  wire n6589;
  wire n6592;
  wire n6595;
  wire n6598;
  wire n6601;
  wire n6604;
  wire n6607;
  wire n6610;
  wire n6613;
  wire n6616;
  wire n6619;
  wire n6622;
  wire n6625;
  wire n6628;
  wire n6631;
  wire n6634;
  wire n6637;
  wire n6640;
  wire n6643;
  wire n6646;
  wire n6649;
  wire n6652;
  wire [31:0] n6654;
  reg [17:0] n6655;
  assign y = y1; //(module output)
  /* fppow16.vhdl:626:8  */
  assign y0 = n6655; // (signal)
  /* fppow16.vhdl:628:8  */
  assign y1 = y0; // (signal)
  /* fppow16.vhdl:632:28  */
  assign n6559 = x == 5'b00000;
  /* fppow16.vhdl:633:28  */
  assign n6562 = x == 5'b00001;
  /* fppow16.vhdl:634:28  */
  assign n6565 = x == 5'b00010;
  /* fppow16.vhdl:635:28  */
  assign n6568 = x == 5'b00011;
  /* fppow16.vhdl:636:28  */
  assign n6571 = x == 5'b00100;
  /* fppow16.vhdl:637:28  */
  assign n6574 = x == 5'b00101;
  /* fppow16.vhdl:638:28  */
  assign n6577 = x == 5'b00110;
  /* fppow16.vhdl:639:28  */
  assign n6580 = x == 5'b00111;
  /* fppow16.vhdl:640:28  */
  assign n6583 = x == 5'b01000;
  /* fppow16.vhdl:641:28  */
  assign n6586 = x == 5'b01001;
  /* fppow16.vhdl:642:28  */
  assign n6589 = x == 5'b01010;
  /* fppow16.vhdl:643:28  */
  assign n6592 = x == 5'b01011;
  /* fppow16.vhdl:644:28  */
  assign n6595 = x == 5'b01100;
  /* fppow16.vhdl:645:28  */
  assign n6598 = x == 5'b01101;
  /* fppow16.vhdl:646:28  */
  assign n6601 = x == 5'b01110;
  /* fppow16.vhdl:647:28  */
  assign n6604 = x == 5'b01111;
  /* fppow16.vhdl:648:28  */
  assign n6607 = x == 5'b10000;
  /* fppow16.vhdl:649:28  */
  assign n6610 = x == 5'b10001;
  /* fppow16.vhdl:650:28  */
  assign n6613 = x == 5'b10010;
  /* fppow16.vhdl:651:28  */
  assign n6616 = x == 5'b10011;
  /* fppow16.vhdl:652:28  */
  assign n6619 = x == 5'b10100;
  /* fppow16.vhdl:653:28  */
  assign n6622 = x == 5'b10101;
  /* fppow16.vhdl:654:28  */
  assign n6625 = x == 5'b10110;
  /* fppow16.vhdl:655:28  */
  assign n6628 = x == 5'b10111;
  /* fppow16.vhdl:656:28  */
  assign n6631 = x == 5'b11000;
  /* fppow16.vhdl:657:28  */
  assign n6634 = x == 5'b11001;
  /* fppow16.vhdl:658:28  */
  assign n6637 = x == 5'b11010;
  /* fppow16.vhdl:659:28  */
  assign n6640 = x == 5'b11011;
  /* fppow16.vhdl:660:28  */
  assign n6643 = x == 5'b11100;
  /* fppow16.vhdl:661:28  */
  assign n6646 = x == 5'b11101;
  /* fppow16.vhdl:662:28  */
  assign n6649 = x == 5'b11110;
  /* fppow16.vhdl:663:28  */
  assign n6652 = x == 5'b11111;
  assign n6654 = {n6652, n6649, n6646, n6643, n6640, n6637, n6634, n6631, n6628, n6625, n6622, n6619, n6616, n6613, n6610, n6607, n6604, n6601, n6598, n6595, n6592, n6589, n6586, n6583, n6580, n6577, n6574, n6571, n6568, n6565, n6562, n6559};
  /* fppow16.vhdl:631:4  */
  always @*
    case (n6654)
      32'b10000000000000000000000000000000: n6655 = 18'b101010111110011010;
      32'b01000000000000000000000000000000: n6655 = 18'b101001100101101100;
      32'b00100000000000000000000000000000: n6655 = 18'b101000001100111110;
      32'b00010000000000000000000000000000: n6655 = 18'b100110110100001111;
      32'b00001000000000000000000000000000: n6655 = 18'b100101011011100001;
      32'b00000100000000000000000000000000: n6655 = 18'b100100000010110011;
      32'b00000010000000000000000000000000: n6655 = 18'b100010101010000101;
      32'b00000001000000000000000000000000: n6655 = 18'b100001010001010110;
      32'b00000000100000000000000000000000: n6655 = 18'b011111111000101000;
      32'b00000000010000000000000000000000: n6655 = 18'b011110011111111010;
      32'b00000000001000000000000000000000: n6655 = 18'b011101000111001011;
      32'b00000000000100000000000000000000: n6655 = 18'b011011101110011101;
      32'b00000000000010000000000000000000: n6655 = 18'b011010010101101111;
      32'b00000000000001000000000000000000: n6655 = 18'b011000111101000001;
      32'b00000000000000100000000000000000: n6655 = 18'b010111100100010010;
      32'b00000000000000010000000000000000: n6655 = 18'b010110001011100100;
      32'b00000000000000001000000000000000: n6655 = 18'b010100110010110110;
      32'b00000000000000000100000000000000: n6655 = 18'b010011011010001000;
      32'b00000000000000000010000000000000: n6655 = 18'b010010000001011001;
      32'b00000000000000000001000000000000: n6655 = 18'b010000101000101011;
      32'b00000000000000000000100000000000: n6655 = 18'b001111001111111101;
      32'b00000000000000000000010000000000: n6655 = 18'b001101110111001111;
      32'b00000000000000000000001000000000: n6655 = 18'b001100011110100000;
      32'b00000000000000000000000100000000: n6655 = 18'b001011000101110010;
      32'b00000000000000000000000010000000: n6655 = 18'b001001101101000100;
      32'b00000000000000000000000001000000: n6655 = 18'b001000010100010110;
      32'b00000000000000000000000000100000: n6655 = 18'b000110111011100111;
      32'b00000000000000000000000000010000: n6655 = 18'b000101100010111001;
      32'b00000000000000000000000000001000: n6655 = 18'b000100001010001011;
      32'b00000000000000000000000000000100: n6655 = 18'b000010110001011101;
      32'b00000000000000000000000000000010: n6655 = 18'b000001011000101110;
      32'b00000000000000000000000000000001: n6655 = 18'b000000000000000000;
      default: n6655 = 18'bX;
    endcase
endmodule

module intadder_9_freq500_uid82
  (input  clk,
   input  [8:0] x,
   input  [8:0] y,
   input  cin,
   output [8:0] r);
  wire [8:0] rtmp;
  wire [8:0] x_d1;
  wire [8:0] y_d1;
  wire cin_d1;
  wire cin_d2;
  wire cin_d3;
  wire cin_d4;
  wire cin_d5;
  wire cin_d6;
  wire cin_d7;
  wire cin_d8;
  wire cin_d9;
  wire cin_d10;
  wire cin_d11;
  wire cin_d12;
  wire cin_d13;
  wire cin_d14;
  wire cin_d15;
  wire [8:0] n6536;
  wire [8:0] n6537;
  wire [8:0] n6538;
  reg [8:0] n6539;
  reg [8:0] n6540;
  reg n6541;
  reg n6542;
  reg n6543;
  reg n6544;
  reg n6545;
  reg n6546;
  reg n6547;
  reg n6548;
  reg n6549;
  reg n6550;
  reg n6551;
  reg n6552;
  reg n6553;
  reg n6554;
  reg n6555;
  assign r = rtmp; //(module output)
  /* fppow16.vhdl:3784:8  */
  assign rtmp = n6538; // (signal)
  /* fppow16.vhdl:3786:8  */
  assign x_d1 = n6539; // (signal)
  /* fppow16.vhdl:3788:8  */
  assign y_d1 = n6540; // (signal)
  /* fppow16.vhdl:3790:8  */
  assign cin_d1 = n6541; // (signal)
  /* fppow16.vhdl:3790:16  */
  assign cin_d2 = n6542; // (signal)
  /* fppow16.vhdl:3790:24  */
  assign cin_d3 = n6543; // (signal)
  /* fppow16.vhdl:3790:32  */
  assign cin_d4 = n6544; // (signal)
  /* fppow16.vhdl:3790:40  */
  assign cin_d5 = n6545; // (signal)
  /* fppow16.vhdl:3790:48  */
  assign cin_d6 = n6546; // (signal)
  /* fppow16.vhdl:3790:56  */
  assign cin_d7 = n6547; // (signal)
  /* fppow16.vhdl:3790:64  */
  assign cin_d8 = n6548; // (signal)
  /* fppow16.vhdl:3790:72  */
  assign cin_d9 = n6549; // (signal)
  /* fppow16.vhdl:3790:80  */
  assign cin_d10 = n6550; // (signal)
  /* fppow16.vhdl:3790:89  */
  assign cin_d11 = n6551; // (signal)
  /* fppow16.vhdl:3790:98  */
  assign cin_d12 = n6552; // (signal)
  /* fppow16.vhdl:3790:107  */
  assign cin_d13 = n6553; // (signal)
  /* fppow16.vhdl:3790:116  */
  assign cin_d14 = n6554; // (signal)
  /* fppow16.vhdl:3790:125  */
  assign cin_d15 = n6555; // (signal)
  /* fppow16.vhdl:3815:17  */
  assign n6536 = x_d1 + y_d1;
  /* fppow16.vhdl:3815:24  */
  assign n6537 = {8'b0, cin_d15};  //  uext
  /* fppow16.vhdl:3815:24  */
  assign n6538 = n6536 + n6537;
  /* fppow16.vhdl:3795:10  */
  always @(posedge clk)
    n6539 <= x;
  /* fppow16.vhdl:3795:10  */
  always @(posedge clk)
    n6540 <= y;
  /* fppow16.vhdl:3795:10  */
  always @(posedge clk)
    n6541 <= cin;
  /* fppow16.vhdl:3795:10  */
  always @(posedge clk)
    n6542 <= cin_d1;
  /* fppow16.vhdl:3795:10  */
  always @(posedge clk)
    n6543 <= cin_d2;
  /* fppow16.vhdl:3795:10  */
  always @(posedge clk)
    n6544 <= cin_d3;
  /* fppow16.vhdl:3795:10  */
  always @(posedge clk)
    n6545 <= cin_d4;
  /* fppow16.vhdl:3795:10  */
  always @(posedge clk)
    n6546 <= cin_d5;
  /* fppow16.vhdl:3795:10  */
  always @(posedge clk)
    n6547 <= cin_d6;
  /* fppow16.vhdl:3795:10  */
  always @(posedge clk)
    n6548 <= cin_d7;
  /* fppow16.vhdl:3795:10  */
  always @(posedge clk)
    n6549 <= cin_d8;
  /* fppow16.vhdl:3795:10  */
  always @(posedge clk)
    n6550 <= cin_d9;
  /* fppow16.vhdl:3795:10  */
  always @(posedge clk)
    n6551 <= cin_d10;
  /* fppow16.vhdl:3795:10  */
  always @(posedge clk)
    n6552 <= cin_d11;
  /* fppow16.vhdl:3795:10  */
  always @(posedge clk)
    n6553 <= cin_d12;
  /* fppow16.vhdl:3795:10  */
  always @(posedge clk)
    n6554 <= cin_d13;
  /* fppow16.vhdl:3795:10  */
  always @(posedge clk)
    n6555 <= cin_d14;
endmodule

module fixrealkcm_freq500_uid72_t1_freq500_uid78
  (input  [1:0] x,
   output [3:0] y);
  wire [3:0] y0;
  wire [3:0] y1;
  wire n6501;
  wire n6504;
  wire n6507;
  wire n6510;
  wire [3:0] n6512;
  reg [3:0] n6513;
  assign y = y1; //(module output)
  /* fppow16.vhdl:582:8  */
  assign y0 = n6513; // (signal)
  /* fppow16.vhdl:584:8  */
  assign y1 = y0; // (signal)
  /* fppow16.vhdl:588:14  */
  assign n6501 = x == 2'b00;
  /* fppow16.vhdl:589:14  */
  assign n6504 = x == 2'b01;
  /* fppow16.vhdl:590:14  */
  assign n6507 = x == 2'b10;
  /* fppow16.vhdl:591:14  */
  assign n6510 = x == 2'b11;
  assign n6512 = {n6510, n6507, n6504, n6501};
  /* fppow16.vhdl:587:4  */
  always @*
    case (n6512)
      4'b1000: n6513 = 4'b1001;
      4'b0100: n6513 = 4'b0110;
      4'b0010: n6513 = 4'b0011;
      4'b0001: n6513 = 4'b0000;
      default: n6513 = 4'bX;
    endcase
endmodule

module fixrealkcm_freq500_uid72_t0_freq500_uid75
  (input  [4:0] x,
   output [8:0] y);
  wire [8:0] y0;
  wire [8:0] y1;
  wire n6401;
  wire n6404;
  wire n6407;
  wire n6410;
  wire n6413;
  wire n6416;
  wire n6419;
  wire n6422;
  wire n6425;
  wire n6428;
  wire n6431;
  wire n6434;
  wire n6437;
  wire n6440;
  wire n6443;
  wire n6446;
  wire n6449;
  wire n6452;
  wire n6455;
  wire n6458;
  wire n6461;
  wire n6464;
  wire n6467;
  wire n6470;
  wire n6473;
  wire n6476;
  wire n6479;
  wire n6482;
  wire n6485;
  wire n6488;
  wire n6491;
  wire n6494;
  wire [31:0] n6496;
  reg [8:0] n6497;
  assign y = y1; //(module output)
  /* fppow16.vhdl:510:8  */
  assign y0 = n6497; // (signal)
  /* fppow16.vhdl:512:8  */
  assign y1 = y0; // (signal)
  /* fppow16.vhdl:516:19  */
  assign n6401 = x == 5'b00000;
  /* fppow16.vhdl:517:19  */
  assign n6404 = x == 5'b00001;
  /* fppow16.vhdl:518:19  */
  assign n6407 = x == 5'b00010;
  /* fppow16.vhdl:519:19  */
  assign n6410 = x == 5'b00011;
  /* fppow16.vhdl:520:19  */
  assign n6413 = x == 5'b00100;
  /* fppow16.vhdl:521:19  */
  assign n6416 = x == 5'b00101;
  /* fppow16.vhdl:522:19  */
  assign n6419 = x == 5'b00110;
  /* fppow16.vhdl:523:19  */
  assign n6422 = x == 5'b00111;
  /* fppow16.vhdl:524:19  */
  assign n6425 = x == 5'b01000;
  /* fppow16.vhdl:525:19  */
  assign n6428 = x == 5'b01001;
  /* fppow16.vhdl:526:19  */
  assign n6431 = x == 5'b01010;
  /* fppow16.vhdl:527:19  */
  assign n6434 = x == 5'b01011;
  /* fppow16.vhdl:528:19  */
  assign n6437 = x == 5'b01100;
  /* fppow16.vhdl:529:19  */
  assign n6440 = x == 5'b01101;
  /* fppow16.vhdl:530:19  */
  assign n6443 = x == 5'b01110;
  /* fppow16.vhdl:531:19  */
  assign n6446 = x == 5'b01111;
  /* fppow16.vhdl:532:19  */
  assign n6449 = x == 5'b10000;
  /* fppow16.vhdl:533:19  */
  assign n6452 = x == 5'b10001;
  /* fppow16.vhdl:534:19  */
  assign n6455 = x == 5'b10010;
  /* fppow16.vhdl:535:19  */
  assign n6458 = x == 5'b10011;
  /* fppow16.vhdl:536:19  */
  assign n6461 = x == 5'b10100;
  /* fppow16.vhdl:537:19  */
  assign n6464 = x == 5'b10101;
  /* fppow16.vhdl:538:19  */
  assign n6467 = x == 5'b10110;
  /* fppow16.vhdl:539:19  */
  assign n6470 = x == 5'b10111;
  /* fppow16.vhdl:540:19  */
  assign n6473 = x == 5'b11000;
  /* fppow16.vhdl:541:19  */
  assign n6476 = x == 5'b11001;
  /* fppow16.vhdl:542:19  */
  assign n6479 = x == 5'b11010;
  /* fppow16.vhdl:543:19  */
  assign n6482 = x == 5'b11011;
  /* fppow16.vhdl:544:19  */
  assign n6485 = x == 5'b11100;
  /* fppow16.vhdl:545:19  */
  assign n6488 = x == 5'b11101;
  /* fppow16.vhdl:546:19  */
  assign n6491 = x == 5'b11110;
  /* fppow16.vhdl:547:19  */
  assign n6494 = x == 5'b11111;
  assign n6496 = {n6494, n6491, n6488, n6485, n6482, n6479, n6476, n6473, n6470, n6467, n6464, n6461, n6458, n6455, n6452, n6449, n6446, n6443, n6440, n6437, n6434, n6431, n6428, n6425, n6422, n6419, n6416, n6413, n6410, n6407, n6404, n6401};
  /* fppow16.vhdl:515:4  */
  always @*
    case (n6496)
      32'b10000000000000000000000000000000: n6497 = 9'b101101110;
      32'b01000000000000000000000000000000: n6497 = 9'b101100010;
      32'b00100000000000000000000000000000: n6497 = 9'b101010111;
      32'b00010000000000000000000000000000: n6497 = 9'b101001011;
      32'b00001000000000000000000000000000: n6497 = 9'b101000000;
      32'b00000100000000000000000000000000: n6497 = 9'b100110100;
      32'b00000010000000000000000000000000: n6497 = 9'b100101001;
      32'b00000001000000000000000000000000: n6497 = 9'b100011101;
      32'b00000000100000000000000000000000: n6497 = 9'b100010001;
      32'b00000000010000000000000000000000: n6497 = 9'b100000110;
      32'b00000000001000000000000000000000: n6497 = 9'b011111010;
      32'b00000000000100000000000000000000: n6497 = 9'b011101111;
      32'b00000000000010000000000000000000: n6497 = 9'b011100011;
      32'b00000000000001000000000000000000: n6497 = 9'b011011000;
      32'b00000000000000100000000000000000: n6497 = 9'b011001100;
      32'b00000000000000010000000000000000: n6497 = 9'b011000001;
      32'b00000000000000001000000000000000: n6497 = 9'b010110101;
      32'b00000000000000000100000000000000: n6497 = 9'b010101010;
      32'b00000000000000000010000000000000: n6497 = 9'b010011110;
      32'b00000000000000000001000000000000: n6497 = 9'b010010010;
      32'b00000000000000000000100000000000: n6497 = 9'b010000111;
      32'b00000000000000000000010000000000: n6497 = 9'b001111011;
      32'b00000000000000000000001000000000: n6497 = 9'b001110000;
      32'b00000000000000000000000100000000: n6497 = 9'b001100100;
      32'b00000000000000000000000010000000: n6497 = 9'b001011001;
      32'b00000000000000000000000001000000: n6497 = 9'b001001101;
      32'b00000000000000000000000000100000: n6497 = 9'b001000010;
      32'b00000000000000000000000000010000: n6497 = 9'b000110110;
      32'b00000000000000000000000000001000: n6497 = 9'b000101011;
      32'b00000000000000000000000000000100: n6497 = 9'b000011111;
      32'b00000000000000000000000000000010: n6497 = 9'b000010100;
      32'b00000000000000000000000000000001: n6497 = 9'b000001000;
      default: n6497 = 9'bX;
    endcase
endmodule

module intadder_14_freq500_uid108
  (input  clk,
   input  [13:0] x,
   input  [13:0] y,
   input  cin,
   output [13:0] r);
  wire [13:0] rtmp;
  wire [13:0] x_d1;
  wire [13:0] y_d1;
  wire cin_d1;
  wire cin_d2;
  wire cin_d3;
  wire cin_d4;
  wire cin_d5;
  wire cin_d6;
  wire cin_d7;
  wire cin_d8;
  wire cin_d9;
  wire cin_d10;
  wire cin_d11;
  wire cin_d12;
  wire cin_d13;
  wire cin_d14;
  wire cin_d15;
  wire cin_d16;
  wire cin_d17;
  wire [13:0] n6376;
  wire [13:0] n6377;
  wire [13:0] n6378;
  reg [13:0] n6379;
  reg [13:0] n6380;
  reg n6381;
  reg n6382;
  reg n6383;
  reg n6384;
  reg n6385;
  reg n6386;
  reg n6387;
  reg n6388;
  reg n6389;
  reg n6390;
  reg n6391;
  reg n6392;
  reg n6393;
  reg n6394;
  reg n6395;
  reg n6396;
  reg n6397;
  assign r = rtmp; //(module output)
  /* fppow16.vhdl:4310:8  */
  assign rtmp = n6378; // (signal)
  /* fppow16.vhdl:4312:8  */
  assign x_d1 = n6379; // (signal)
  /* fppow16.vhdl:4314:8  */
  assign y_d1 = n6380; // (signal)
  /* fppow16.vhdl:4316:8  */
  assign cin_d1 = n6381; // (signal)
  /* fppow16.vhdl:4316:16  */
  assign cin_d2 = n6382; // (signal)
  /* fppow16.vhdl:4316:24  */
  assign cin_d3 = n6383; // (signal)
  /* fppow16.vhdl:4316:32  */
  assign cin_d4 = n6384; // (signal)
  /* fppow16.vhdl:4316:40  */
  assign cin_d5 = n6385; // (signal)
  /* fppow16.vhdl:4316:48  */
  assign cin_d6 = n6386; // (signal)
  /* fppow16.vhdl:4316:56  */
  assign cin_d7 = n6387; // (signal)
  /* fppow16.vhdl:4316:64  */
  assign cin_d8 = n6388; // (signal)
  /* fppow16.vhdl:4316:72  */
  assign cin_d9 = n6389; // (signal)
  /* fppow16.vhdl:4316:80  */
  assign cin_d10 = n6390; // (signal)
  /* fppow16.vhdl:4316:89  */
  assign cin_d11 = n6391; // (signal)
  /* fppow16.vhdl:4316:98  */
  assign cin_d12 = n6392; // (signal)
  /* fppow16.vhdl:4316:107  */
  assign cin_d13 = n6393; // (signal)
  /* fppow16.vhdl:4316:116  */
  assign cin_d14 = n6394; // (signal)
  /* fppow16.vhdl:4316:125  */
  assign cin_d15 = n6395; // (signal)
  /* fppow16.vhdl:4316:134  */
  assign cin_d16 = n6396; // (signal)
  /* fppow16.vhdl:4316:143  */
  assign cin_d17 = n6397; // (signal)
  /* fppow16.vhdl:4343:17  */
  assign n6376 = x_d1 + y_d1;
  /* fppow16.vhdl:4343:24  */
  assign n6377 = {13'b0, cin_d17};  //  uext
  /* fppow16.vhdl:4343:24  */
  assign n6378 = n6376 + n6377;
  /* fppow16.vhdl:4321:10  */
  always @(posedge clk)
    n6379 <= x;
  /* fppow16.vhdl:4321:10  */
  always @(posedge clk)
    n6380 <= y;
  /* fppow16.vhdl:4321:10  */
  always @(posedge clk)
    n6381 <= cin;
  /* fppow16.vhdl:4321:10  */
  always @(posedge clk)
    n6382 <= cin_d1;
  /* fppow16.vhdl:4321:10  */
  always @(posedge clk)
    n6383 <= cin_d2;
  /* fppow16.vhdl:4321:10  */
  always @(posedge clk)
    n6384 <= cin_d3;
  /* fppow16.vhdl:4321:10  */
  always @(posedge clk)
    n6385 <= cin_d4;
  /* fppow16.vhdl:4321:10  */
  always @(posedge clk)
    n6386 <= cin_d5;
  /* fppow16.vhdl:4321:10  */
  always @(posedge clk)
    n6387 <= cin_d6;
  /* fppow16.vhdl:4321:10  */
  always @(posedge clk)
    n6388 <= cin_d7;
  /* fppow16.vhdl:4321:10  */
  always @(posedge clk)
    n6389 <= cin_d8;
  /* fppow16.vhdl:4321:10  */
  always @(posedge clk)
    n6390 <= cin_d9;
  /* fppow16.vhdl:4321:10  */
  always @(posedge clk)
    n6391 <= cin_d10;
  /* fppow16.vhdl:4321:10  */
  always @(posedge clk)
    n6392 <= cin_d11;
  /* fppow16.vhdl:4321:10  */
  always @(posedge clk)
    n6393 <= cin_d12;
  /* fppow16.vhdl:4321:10  */
  always @(posedge clk)
    n6394 <= cin_d13;
  /* fppow16.vhdl:4321:10  */
  always @(posedge clk)
    n6395 <= cin_d14;
  /* fppow16.vhdl:4321:10  */
  always @(posedge clk)
    n6396 <= cin_d15;
  /* fppow16.vhdl:4321:10  */
  always @(posedge clk)
    n6397 <= cin_d16;
endmodule

module intmultiplier_3x4_5_freq500_uid104
  (input  clk,
   input  [2:0] x,
   input  [3:0] y,
   output [4:0] r);
  wire [2:0] xx;
  wire [3:0] yy;
  wire [6:0] rr;
  wire [6:0] n6348;
  wire [6:0] n6349;
  wire [6:0] n6350;
  wire [4:0] n6351;
  assign r = n6351; //(module output)
  /* fppow16.vhdl:4267:8  */
  assign rr = n6350; // (signal)
  /* fppow16.vhdl:4274:12  */
  assign n6348 = {4'b0, xx};  //  uext
  /* fppow16.vhdl:4274:12  */
  assign n6349 = {3'b0, yy};  //  uext
  /* fppow16.vhdl:4274:12  */
  assign n6350 = n6348 * n6349; // umul
  /* fppow16.vhdl:4275:28  */
  assign n6351 = rr[6:2]; // extract
endmodule

module intadder_4_freq500_uid102
  (input  clk,
   input  [3:0] x,
   input  [3:0] y,
   input  cin,
   output [3:0] r);
  wire [3:0] rtmp;
  wire [3:0] y_d1;
  wire [3:0] y_d2;
  wire [3:0] y_d3;
  wire [3:0] y_d4;
  wire [3:0] y_d5;
  wire [3:0] y_d6;
  wire [3:0] y_d7;
  wire [3:0] y_d8;
  wire [3:0] y_d9;
  wire [3:0] y_d10;
  wire [3:0] y_d11;
  wire [3:0] y_d12;
  wire [3:0] y_d13;
  wire [3:0] y_d14;
  wire [3:0] y_d15;
  wire [3:0] y_d16;
  wire cin_d1;
  wire cin_d2;
  wire cin_d3;
  wire cin_d4;
  wire cin_d5;
  wire cin_d6;
  wire cin_d7;
  wire cin_d8;
  wire cin_d9;
  wire cin_d10;
  wire cin_d11;
  wire cin_d12;
  wire cin_d13;
  wire cin_d14;
  wire cin_d15;
  wire cin_d16;
  wire [3:0] n6312;
  wire [3:0] n6313;
  wire [3:0] n6314;
  reg [3:0] n6315;
  reg [3:0] n6316;
  reg [3:0] n6317;
  reg [3:0] n6318;
  reg [3:0] n6319;
  reg [3:0] n6320;
  reg [3:0] n6321;
  reg [3:0] n6322;
  reg [3:0] n6323;
  reg [3:0] n6324;
  reg [3:0] n6325;
  reg [3:0] n6326;
  reg [3:0] n6327;
  reg [3:0] n6328;
  reg [3:0] n6329;
  reg [3:0] n6330;
  reg n6331;
  reg n6332;
  reg n6333;
  reg n6334;
  reg n6335;
  reg n6336;
  reg n6337;
  reg n6338;
  reg n6339;
  reg n6340;
  reg n6341;
  reg n6342;
  reg n6343;
  reg n6344;
  reg n6345;
  reg n6346;
  assign r = rtmp; //(module output)
  /* fppow16.vhdl:4181:8  */
  assign rtmp = n6314; // (signal)
  /* fppow16.vhdl:4183:8  */
  assign y_d1 = n6315; // (signal)
  /* fppow16.vhdl:4183:14  */
  assign y_d2 = n6316; // (signal)
  /* fppow16.vhdl:4183:20  */
  assign y_d3 = n6317; // (signal)
  /* fppow16.vhdl:4183:26  */
  assign y_d4 = n6318; // (signal)
  /* fppow16.vhdl:4183:32  */
  assign y_d5 = n6319; // (signal)
  /* fppow16.vhdl:4183:38  */
  assign y_d6 = n6320; // (signal)
  /* fppow16.vhdl:4183:44  */
  assign y_d7 = n6321; // (signal)
  /* fppow16.vhdl:4183:50  */
  assign y_d8 = n6322; // (signal)
  /* fppow16.vhdl:4183:56  */
  assign y_d9 = n6323; // (signal)
  /* fppow16.vhdl:4183:62  */
  assign y_d10 = n6324; // (signal)
  /* fppow16.vhdl:4183:69  */
  assign y_d11 = n6325; // (signal)
  /* fppow16.vhdl:4183:76  */
  assign y_d12 = n6326; // (signal)
  /* fppow16.vhdl:4183:83  */
  assign y_d13 = n6327; // (signal)
  /* fppow16.vhdl:4183:90  */
  assign y_d14 = n6328; // (signal)
  /* fppow16.vhdl:4183:97  */
  assign y_d15 = n6329; // (signal)
  /* fppow16.vhdl:4183:104  */
  assign y_d16 = n6330; // (signal)
  /* fppow16.vhdl:4185:8  */
  assign cin_d1 = n6331; // (signal)
  /* fppow16.vhdl:4185:16  */
  assign cin_d2 = n6332; // (signal)
  /* fppow16.vhdl:4185:24  */
  assign cin_d3 = n6333; // (signal)
  /* fppow16.vhdl:4185:32  */
  assign cin_d4 = n6334; // (signal)
  /* fppow16.vhdl:4185:40  */
  assign cin_d5 = n6335; // (signal)
  /* fppow16.vhdl:4185:48  */
  assign cin_d6 = n6336; // (signal)
  /* fppow16.vhdl:4185:56  */
  assign cin_d7 = n6337; // (signal)
  /* fppow16.vhdl:4185:64  */
  assign cin_d8 = n6338; // (signal)
  /* fppow16.vhdl:4185:72  */
  assign cin_d9 = n6339; // (signal)
  /* fppow16.vhdl:4185:80  */
  assign cin_d10 = n6340; // (signal)
  /* fppow16.vhdl:4185:89  */
  assign cin_d11 = n6341; // (signal)
  /* fppow16.vhdl:4185:98  */
  assign cin_d12 = n6342; // (signal)
  /* fppow16.vhdl:4185:107  */
  assign cin_d13 = n6343; // (signal)
  /* fppow16.vhdl:4185:116  */
  assign cin_d14 = n6344; // (signal)
  /* fppow16.vhdl:4185:125  */
  assign cin_d15 = n6345; // (signal)
  /* fppow16.vhdl:4185:134  */
  assign cin_d16 = n6346; // (signal)
  /* fppow16.vhdl:4225:14  */
  assign n6312 = x + y_d16;
  /* fppow16.vhdl:4225:22  */
  assign n6313 = {3'b0, cin_d16};  //  uext
  /* fppow16.vhdl:4225:22  */
  assign n6314 = n6312 + n6313;
  /* fppow16.vhdl:4190:10  */
  always @(posedge clk)
    n6315 <= y;
  /* fppow16.vhdl:4190:10  */
  always @(posedge clk)
    n6316 <= y_d1;
  /* fppow16.vhdl:4190:10  */
  always @(posedge clk)
    n6317 <= y_d2;
  /* fppow16.vhdl:4190:10  */
  always @(posedge clk)
    n6318 <= y_d3;
  /* fppow16.vhdl:4190:10  */
  always @(posedge clk)
    n6319 <= y_d4;
  /* fppow16.vhdl:4190:10  */
  always @(posedge clk)
    n6320 <= y_d5;
  /* fppow16.vhdl:4190:10  */
  always @(posedge clk)
    n6321 <= y_d6;
  /* fppow16.vhdl:4190:10  */
  always @(posedge clk)
    n6322 <= y_d7;
  /* fppow16.vhdl:4190:10  */
  always @(posedge clk)
    n6323 <= y_d8;
  /* fppow16.vhdl:4190:10  */
  always @(posedge clk)
    n6324 <= y_d9;
  /* fppow16.vhdl:4190:10  */
  always @(posedge clk)
    n6325 <= y_d10;
  /* fppow16.vhdl:4190:10  */
  always @(posedge clk)
    n6326 <= y_d11;
  /* fppow16.vhdl:4190:10  */
  always @(posedge clk)
    n6327 <= y_d12;
  /* fppow16.vhdl:4190:10  */
  always @(posedge clk)
    n6328 <= y_d13;
  /* fppow16.vhdl:4190:10  */
  always @(posedge clk)
    n6329 <= y_d14;
  /* fppow16.vhdl:4190:10  */
  always @(posedge clk)
    n6330 <= y_d15;
  /* fppow16.vhdl:4190:10  */
  always @(posedge clk)
    n6331 <= cin;
  /* fppow16.vhdl:4190:10  */
  always @(posedge clk)
    n6332 <= cin_d1;
  /* fppow16.vhdl:4190:10  */
  always @(posedge clk)
    n6333 <= cin_d2;
  /* fppow16.vhdl:4190:10  */
  always @(posedge clk)
    n6334 <= cin_d3;
  /* fppow16.vhdl:4190:10  */
  always @(posedge clk)
    n6335 <= cin_d4;
  /* fppow16.vhdl:4190:10  */
  always @(posedge clk)
    n6336 <= cin_d5;
  /* fppow16.vhdl:4190:10  */
  always @(posedge clk)
    n6337 <= cin_d6;
  /* fppow16.vhdl:4190:10  */
  always @(posedge clk)
    n6338 <= cin_d7;
  /* fppow16.vhdl:4190:10  */
  always @(posedge clk)
    n6339 <= cin_d8;
  /* fppow16.vhdl:4190:10  */
  always @(posedge clk)
    n6340 <= cin_d9;
  /* fppow16.vhdl:4190:10  */
  always @(posedge clk)
    n6341 <= cin_d10;
  /* fppow16.vhdl:4190:10  */
  always @(posedge clk)
    n6342 <= cin_d11;
  /* fppow16.vhdl:4190:10  */
  always @(posedge clk)
    n6343 <= cin_d12;
  /* fppow16.vhdl:4190:10  */
  always @(posedge clk)
    n6344 <= cin_d13;
  /* fppow16.vhdl:4190:10  */
  always @(posedge clk)
    n6345 <= cin_d14;
  /* fppow16.vhdl:4190:10  */
  always @(posedge clk)
    n6346 <= cin_d15;
endmodule

module fixfunctionbytable_freq500_uid97
  (input  [2:0] x,
   output [2:0] y);
  wire [2:0] y0;
  wire [2:0] y1;
  wire n6250;
  wire n6253;
  wire n6256;
  wire n6259;
  wire n6262;
  wire n6265;
  wire n6268;
  wire n6271;
  wire [7:0] n6273;
  reg [2:0] n6274;
  assign y = y1; //(module output)
  /* fppow16.vhdl:1766:8  */
  assign y0 = n6274; // (signal)
  /* fppow16.vhdl:1768:8  */
  assign y1 = y0; // (signal)
  /* fppow16.vhdl:1772:13  */
  assign n6250 = x == 3'b000;
  /* fppow16.vhdl:1773:13  */
  assign n6253 = x == 3'b001;
  /* fppow16.vhdl:1774:13  */
  assign n6256 = x == 3'b010;
  /* fppow16.vhdl:1775:13  */
  assign n6259 = x == 3'b011;
  /* fppow16.vhdl:1776:13  */
  assign n6262 = x == 3'b100;
  /* fppow16.vhdl:1777:13  */
  assign n6265 = x == 3'b101;
  /* fppow16.vhdl:1778:13  */
  assign n6268 = x == 3'b110;
  /* fppow16.vhdl:1779:13  */
  assign n6271 = x == 3'b111;
  assign n6273 = {n6271, n6268, n6265, n6262, n6259, n6256, n6253, n6250};
  /* fppow16.vhdl:1771:4  */
  always @*
    case (n6273)
      8'b10000000: n6274 = 3'b111;
      8'b01000000: n6274 = 3'b110;
      8'b00100000: n6274 = 3'b101;
      8'b00010000: n6274 = 3'b100;
      8'b00001000: n6274 = 3'b011;
      8'b00000100: n6274 = 3'b010;
      8'b00000010: n6274 = 3'b001;
      8'b00000001: n6274 = 3'b000;
      default: n6274 = 3'bX;
    endcase
endmodule

module fixfunctionbytable_freq500_uid94
  (input  [9:0] x,
   output [13:0] y);
  wire [13:0] y0;
  wire [13:0] y1;
  wire n3174;
  wire n3177;
  wire n3180;
  wire n3183;
  wire n3186;
  wire n3189;
  wire n3192;
  wire n3195;
  wire n3198;
  wire n3201;
  wire n3204;
  wire n3207;
  wire n3210;
  wire n3213;
  wire n3216;
  wire n3219;
  wire n3222;
  wire n3225;
  wire n3228;
  wire n3231;
  wire n3234;
  wire n3237;
  wire n3240;
  wire n3243;
  wire n3246;
  wire n3249;
  wire n3252;
  wire n3255;
  wire n3258;
  wire n3261;
  wire n3264;
  wire n3267;
  wire n3270;
  wire n3273;
  wire n3276;
  wire n3279;
  wire n3282;
  wire n3285;
  wire n3288;
  wire n3291;
  wire n3294;
  wire n3297;
  wire n3300;
  wire n3303;
  wire n3306;
  wire n3309;
  wire n3312;
  wire n3315;
  wire n3318;
  wire n3321;
  wire n3324;
  wire n3327;
  wire n3330;
  wire n3333;
  wire n3336;
  wire n3339;
  wire n3342;
  wire n3345;
  wire n3348;
  wire n3351;
  wire n3354;
  wire n3357;
  wire n3360;
  wire n3363;
  wire n3366;
  wire n3369;
  wire n3372;
  wire n3375;
  wire n3378;
  wire n3381;
  wire n3384;
  wire n3387;
  wire n3390;
  wire n3393;
  wire n3396;
  wire n3399;
  wire n3402;
  wire n3405;
  wire n3408;
  wire n3411;
  wire n3414;
  wire n3417;
  wire n3420;
  wire n3423;
  wire n3426;
  wire n3429;
  wire n3432;
  wire n3435;
  wire n3438;
  wire n3441;
  wire n3444;
  wire n3447;
  wire n3450;
  wire n3453;
  wire n3456;
  wire n3459;
  wire n3462;
  wire n3465;
  wire n3468;
  wire n3471;
  wire n3474;
  wire n3477;
  wire n3480;
  wire n3483;
  wire n3486;
  wire n3489;
  wire n3492;
  wire n3495;
  wire n3498;
  wire n3501;
  wire n3504;
  wire n3507;
  wire n3510;
  wire n3513;
  wire n3516;
  wire n3519;
  wire n3522;
  wire n3525;
  wire n3528;
  wire n3531;
  wire n3534;
  wire n3537;
  wire n3540;
  wire n3543;
  wire n3546;
  wire n3549;
  wire n3552;
  wire n3555;
  wire n3558;
  wire n3561;
  wire n3564;
  wire n3567;
  wire n3570;
  wire n3573;
  wire n3576;
  wire n3579;
  wire n3582;
  wire n3585;
  wire n3588;
  wire n3591;
  wire n3594;
  wire n3597;
  wire n3600;
  wire n3603;
  wire n3606;
  wire n3609;
  wire n3612;
  wire n3615;
  wire n3618;
  wire n3621;
  wire n3624;
  wire n3627;
  wire n3630;
  wire n3633;
  wire n3636;
  wire n3639;
  wire n3642;
  wire n3645;
  wire n3648;
  wire n3651;
  wire n3654;
  wire n3657;
  wire n3660;
  wire n3663;
  wire n3666;
  wire n3669;
  wire n3672;
  wire n3675;
  wire n3678;
  wire n3681;
  wire n3684;
  wire n3687;
  wire n3690;
  wire n3693;
  wire n3696;
  wire n3699;
  wire n3702;
  wire n3705;
  wire n3708;
  wire n3711;
  wire n3714;
  wire n3717;
  wire n3720;
  wire n3723;
  wire n3726;
  wire n3729;
  wire n3732;
  wire n3735;
  wire n3738;
  wire n3741;
  wire n3744;
  wire n3747;
  wire n3750;
  wire n3753;
  wire n3756;
  wire n3759;
  wire n3762;
  wire n3765;
  wire n3768;
  wire n3771;
  wire n3774;
  wire n3777;
  wire n3780;
  wire n3783;
  wire n3786;
  wire n3789;
  wire n3792;
  wire n3795;
  wire n3798;
  wire n3801;
  wire n3804;
  wire n3807;
  wire n3810;
  wire n3813;
  wire n3816;
  wire n3819;
  wire n3822;
  wire n3825;
  wire n3828;
  wire n3831;
  wire n3834;
  wire n3837;
  wire n3840;
  wire n3843;
  wire n3846;
  wire n3849;
  wire n3852;
  wire n3855;
  wire n3858;
  wire n3861;
  wire n3864;
  wire n3867;
  wire n3870;
  wire n3873;
  wire n3876;
  wire n3879;
  wire n3882;
  wire n3885;
  wire n3888;
  wire n3891;
  wire n3894;
  wire n3897;
  wire n3900;
  wire n3903;
  wire n3906;
  wire n3909;
  wire n3912;
  wire n3915;
  wire n3918;
  wire n3921;
  wire n3924;
  wire n3927;
  wire n3930;
  wire n3933;
  wire n3936;
  wire n3939;
  wire n3942;
  wire n3945;
  wire n3948;
  wire n3951;
  wire n3954;
  wire n3957;
  wire n3960;
  wire n3963;
  wire n3966;
  wire n3969;
  wire n3972;
  wire n3975;
  wire n3978;
  wire n3981;
  wire n3984;
  wire n3987;
  wire n3990;
  wire n3993;
  wire n3996;
  wire n3999;
  wire n4002;
  wire n4005;
  wire n4008;
  wire n4011;
  wire n4014;
  wire n4017;
  wire n4020;
  wire n4023;
  wire n4026;
  wire n4029;
  wire n4032;
  wire n4035;
  wire n4038;
  wire n4041;
  wire n4044;
  wire n4047;
  wire n4050;
  wire n4053;
  wire n4056;
  wire n4059;
  wire n4062;
  wire n4065;
  wire n4068;
  wire n4071;
  wire n4074;
  wire n4077;
  wire n4080;
  wire n4083;
  wire n4086;
  wire n4089;
  wire n4092;
  wire n4095;
  wire n4098;
  wire n4101;
  wire n4104;
  wire n4107;
  wire n4110;
  wire n4113;
  wire n4116;
  wire n4119;
  wire n4122;
  wire n4125;
  wire n4128;
  wire n4131;
  wire n4134;
  wire n4137;
  wire n4140;
  wire n4143;
  wire n4146;
  wire n4149;
  wire n4152;
  wire n4155;
  wire n4158;
  wire n4161;
  wire n4164;
  wire n4167;
  wire n4170;
  wire n4173;
  wire n4176;
  wire n4179;
  wire n4182;
  wire n4185;
  wire n4188;
  wire n4191;
  wire n4194;
  wire n4197;
  wire n4200;
  wire n4203;
  wire n4206;
  wire n4209;
  wire n4212;
  wire n4215;
  wire n4218;
  wire n4221;
  wire n4224;
  wire n4227;
  wire n4230;
  wire n4233;
  wire n4236;
  wire n4239;
  wire n4242;
  wire n4245;
  wire n4248;
  wire n4251;
  wire n4254;
  wire n4257;
  wire n4260;
  wire n4263;
  wire n4266;
  wire n4269;
  wire n4272;
  wire n4275;
  wire n4278;
  wire n4281;
  wire n4284;
  wire n4287;
  wire n4290;
  wire n4293;
  wire n4296;
  wire n4299;
  wire n4302;
  wire n4305;
  wire n4308;
  wire n4311;
  wire n4314;
  wire n4317;
  wire n4320;
  wire n4323;
  wire n4326;
  wire n4329;
  wire n4332;
  wire n4335;
  wire n4338;
  wire n4341;
  wire n4344;
  wire n4347;
  wire n4350;
  wire n4353;
  wire n4356;
  wire n4359;
  wire n4362;
  wire n4365;
  wire n4368;
  wire n4371;
  wire n4374;
  wire n4377;
  wire n4380;
  wire n4383;
  wire n4386;
  wire n4389;
  wire n4392;
  wire n4395;
  wire n4398;
  wire n4401;
  wire n4404;
  wire n4407;
  wire n4410;
  wire n4413;
  wire n4416;
  wire n4419;
  wire n4422;
  wire n4425;
  wire n4428;
  wire n4431;
  wire n4434;
  wire n4437;
  wire n4440;
  wire n4443;
  wire n4446;
  wire n4449;
  wire n4452;
  wire n4455;
  wire n4458;
  wire n4461;
  wire n4464;
  wire n4467;
  wire n4470;
  wire n4473;
  wire n4476;
  wire n4479;
  wire n4482;
  wire n4485;
  wire n4488;
  wire n4491;
  wire n4494;
  wire n4497;
  wire n4500;
  wire n4503;
  wire n4506;
  wire n4509;
  wire n4512;
  wire n4515;
  wire n4518;
  wire n4521;
  wire n4524;
  wire n4527;
  wire n4530;
  wire n4533;
  wire n4536;
  wire n4539;
  wire n4542;
  wire n4545;
  wire n4548;
  wire n4551;
  wire n4554;
  wire n4557;
  wire n4560;
  wire n4563;
  wire n4566;
  wire n4569;
  wire n4572;
  wire n4575;
  wire n4578;
  wire n4581;
  wire n4584;
  wire n4587;
  wire n4590;
  wire n4593;
  wire n4596;
  wire n4599;
  wire n4602;
  wire n4605;
  wire n4608;
  wire n4611;
  wire n4614;
  wire n4617;
  wire n4620;
  wire n4623;
  wire n4626;
  wire n4629;
  wire n4632;
  wire n4635;
  wire n4638;
  wire n4641;
  wire n4644;
  wire n4647;
  wire n4650;
  wire n4653;
  wire n4656;
  wire n4659;
  wire n4662;
  wire n4665;
  wire n4668;
  wire n4671;
  wire n4674;
  wire n4677;
  wire n4680;
  wire n4683;
  wire n4686;
  wire n4689;
  wire n4692;
  wire n4695;
  wire n4698;
  wire n4701;
  wire n4704;
  wire n4707;
  wire n4710;
  wire n4713;
  wire n4716;
  wire n4719;
  wire n4722;
  wire n4725;
  wire n4728;
  wire n4731;
  wire n4734;
  wire n4737;
  wire n4740;
  wire n4743;
  wire n4746;
  wire n4749;
  wire n4752;
  wire n4755;
  wire n4758;
  wire n4761;
  wire n4764;
  wire n4767;
  wire n4770;
  wire n4773;
  wire n4776;
  wire n4779;
  wire n4782;
  wire n4785;
  wire n4788;
  wire n4791;
  wire n4794;
  wire n4797;
  wire n4800;
  wire n4803;
  wire n4806;
  wire n4809;
  wire n4812;
  wire n4815;
  wire n4818;
  wire n4821;
  wire n4824;
  wire n4827;
  wire n4830;
  wire n4833;
  wire n4836;
  wire n4839;
  wire n4842;
  wire n4845;
  wire n4848;
  wire n4851;
  wire n4854;
  wire n4857;
  wire n4860;
  wire n4863;
  wire n4866;
  wire n4869;
  wire n4872;
  wire n4875;
  wire n4878;
  wire n4881;
  wire n4884;
  wire n4887;
  wire n4890;
  wire n4893;
  wire n4896;
  wire n4899;
  wire n4902;
  wire n4905;
  wire n4908;
  wire n4911;
  wire n4914;
  wire n4917;
  wire n4920;
  wire n4923;
  wire n4926;
  wire n4929;
  wire n4932;
  wire n4935;
  wire n4938;
  wire n4941;
  wire n4944;
  wire n4947;
  wire n4950;
  wire n4953;
  wire n4956;
  wire n4959;
  wire n4962;
  wire n4965;
  wire n4968;
  wire n4971;
  wire n4974;
  wire n4977;
  wire n4980;
  wire n4983;
  wire n4986;
  wire n4989;
  wire n4992;
  wire n4995;
  wire n4998;
  wire n5001;
  wire n5004;
  wire n5007;
  wire n5010;
  wire n5013;
  wire n5016;
  wire n5019;
  wire n5022;
  wire n5025;
  wire n5028;
  wire n5031;
  wire n5034;
  wire n5037;
  wire n5040;
  wire n5043;
  wire n5046;
  wire n5049;
  wire n5052;
  wire n5055;
  wire n5058;
  wire n5061;
  wire n5064;
  wire n5067;
  wire n5070;
  wire n5073;
  wire n5076;
  wire n5079;
  wire n5082;
  wire n5085;
  wire n5088;
  wire n5091;
  wire n5094;
  wire n5097;
  wire n5100;
  wire n5103;
  wire n5106;
  wire n5109;
  wire n5112;
  wire n5115;
  wire n5118;
  wire n5121;
  wire n5124;
  wire n5127;
  wire n5130;
  wire n5133;
  wire n5136;
  wire n5139;
  wire n5142;
  wire n5145;
  wire n5148;
  wire n5151;
  wire n5154;
  wire n5157;
  wire n5160;
  wire n5163;
  wire n5166;
  wire n5169;
  wire n5172;
  wire n5175;
  wire n5178;
  wire n5181;
  wire n5184;
  wire n5187;
  wire n5190;
  wire n5193;
  wire n5196;
  wire n5199;
  wire n5202;
  wire n5205;
  wire n5208;
  wire n5211;
  wire n5214;
  wire n5217;
  wire n5220;
  wire n5223;
  wire n5226;
  wire n5229;
  wire n5232;
  wire n5235;
  wire n5238;
  wire n5241;
  wire n5244;
  wire n5247;
  wire n5250;
  wire n5253;
  wire n5256;
  wire n5259;
  wire n5262;
  wire n5265;
  wire n5268;
  wire n5271;
  wire n5274;
  wire n5277;
  wire n5280;
  wire n5283;
  wire n5286;
  wire n5289;
  wire n5292;
  wire n5295;
  wire n5298;
  wire n5301;
  wire n5304;
  wire n5307;
  wire n5310;
  wire n5313;
  wire n5316;
  wire n5319;
  wire n5322;
  wire n5325;
  wire n5328;
  wire n5331;
  wire n5334;
  wire n5337;
  wire n5340;
  wire n5343;
  wire n5346;
  wire n5349;
  wire n5352;
  wire n5355;
  wire n5358;
  wire n5361;
  wire n5364;
  wire n5367;
  wire n5370;
  wire n5373;
  wire n5376;
  wire n5379;
  wire n5382;
  wire n5385;
  wire n5388;
  wire n5391;
  wire n5394;
  wire n5397;
  wire n5400;
  wire n5403;
  wire n5406;
  wire n5409;
  wire n5412;
  wire n5415;
  wire n5418;
  wire n5421;
  wire n5424;
  wire n5427;
  wire n5430;
  wire n5433;
  wire n5436;
  wire n5439;
  wire n5442;
  wire n5445;
  wire n5448;
  wire n5451;
  wire n5454;
  wire n5457;
  wire n5460;
  wire n5463;
  wire n5466;
  wire n5469;
  wire n5472;
  wire n5475;
  wire n5478;
  wire n5481;
  wire n5484;
  wire n5487;
  wire n5490;
  wire n5493;
  wire n5496;
  wire n5499;
  wire n5502;
  wire n5505;
  wire n5508;
  wire n5511;
  wire n5514;
  wire n5517;
  wire n5520;
  wire n5523;
  wire n5526;
  wire n5529;
  wire n5532;
  wire n5535;
  wire n5538;
  wire n5541;
  wire n5544;
  wire n5547;
  wire n5550;
  wire n5553;
  wire n5556;
  wire n5559;
  wire n5562;
  wire n5565;
  wire n5568;
  wire n5571;
  wire n5574;
  wire n5577;
  wire n5580;
  wire n5583;
  wire n5586;
  wire n5589;
  wire n5592;
  wire n5595;
  wire n5598;
  wire n5601;
  wire n5604;
  wire n5607;
  wire n5610;
  wire n5613;
  wire n5616;
  wire n5619;
  wire n5622;
  wire n5625;
  wire n5628;
  wire n5631;
  wire n5634;
  wire n5637;
  wire n5640;
  wire n5643;
  wire n5646;
  wire n5649;
  wire n5652;
  wire n5655;
  wire n5658;
  wire n5661;
  wire n5664;
  wire n5667;
  wire n5670;
  wire n5673;
  wire n5676;
  wire n5679;
  wire n5682;
  wire n5685;
  wire n5688;
  wire n5691;
  wire n5694;
  wire n5697;
  wire n5700;
  wire n5703;
  wire n5706;
  wire n5709;
  wire n5712;
  wire n5715;
  wire n5718;
  wire n5721;
  wire n5724;
  wire n5727;
  wire n5730;
  wire n5733;
  wire n5736;
  wire n5739;
  wire n5742;
  wire n5745;
  wire n5748;
  wire n5751;
  wire n5754;
  wire n5757;
  wire n5760;
  wire n5763;
  wire n5766;
  wire n5769;
  wire n5772;
  wire n5775;
  wire n5778;
  wire n5781;
  wire n5784;
  wire n5787;
  wire n5790;
  wire n5793;
  wire n5796;
  wire n5799;
  wire n5802;
  wire n5805;
  wire n5808;
  wire n5811;
  wire n5814;
  wire n5817;
  wire n5820;
  wire n5823;
  wire n5826;
  wire n5829;
  wire n5832;
  wire n5835;
  wire n5838;
  wire n5841;
  wire n5844;
  wire n5847;
  wire n5850;
  wire n5853;
  wire n5856;
  wire n5859;
  wire n5862;
  wire n5865;
  wire n5868;
  wire n5871;
  wire n5874;
  wire n5877;
  wire n5880;
  wire n5883;
  wire n5886;
  wire n5889;
  wire n5892;
  wire n5895;
  wire n5898;
  wire n5901;
  wire n5904;
  wire n5907;
  wire n5910;
  wire n5913;
  wire n5916;
  wire n5919;
  wire n5922;
  wire n5925;
  wire n5928;
  wire n5931;
  wire n5934;
  wire n5937;
  wire n5940;
  wire n5943;
  wire n5946;
  wire n5949;
  wire n5952;
  wire n5955;
  wire n5958;
  wire n5961;
  wire n5964;
  wire n5967;
  wire n5970;
  wire n5973;
  wire n5976;
  wire n5979;
  wire n5982;
  wire n5985;
  wire n5988;
  wire n5991;
  wire n5994;
  wire n5997;
  wire n6000;
  wire n6003;
  wire n6006;
  wire n6009;
  wire n6012;
  wire n6015;
  wire n6018;
  wire n6021;
  wire n6024;
  wire n6027;
  wire n6030;
  wire n6033;
  wire n6036;
  wire n6039;
  wire n6042;
  wire n6045;
  wire n6048;
  wire n6051;
  wire n6054;
  wire n6057;
  wire n6060;
  wire n6063;
  wire n6066;
  wire n6069;
  wire n6072;
  wire n6075;
  wire n6078;
  wire n6081;
  wire n6084;
  wire n6087;
  wire n6090;
  wire n6093;
  wire n6096;
  wire n6099;
  wire n6102;
  wire n6105;
  wire n6108;
  wire n6111;
  wire n6114;
  wire n6117;
  wire n6120;
  wire n6123;
  wire n6126;
  wire n6129;
  wire n6132;
  wire n6135;
  wire n6138;
  wire n6141;
  wire n6144;
  wire n6147;
  wire n6150;
  wire n6153;
  wire n6156;
  wire n6159;
  wire n6162;
  wire n6165;
  wire n6168;
  wire n6171;
  wire n6174;
  wire n6177;
  wire n6180;
  wire n6183;
  wire n6186;
  wire n6189;
  wire n6192;
  wire n6195;
  wire n6198;
  wire n6201;
  wire n6204;
  wire n6207;
  wire n6210;
  wire n6213;
  wire n6216;
  wire n6219;
  wire n6222;
  wire n6225;
  wire n6228;
  wire n6231;
  wire n6234;
  wire n6237;
  wire n6240;
  wire n6243;
  wire [1023:0] n6245;
  reg [13:0] n6246;
  assign y = y1; //(module output)
  /* fppow16.vhdl:700:8  */
  assign y0 = n6246; // (signal)
  /* fppow16.vhdl:702:8  */
  assign y1 = y0; // (signal)
  /* fppow16.vhdl:706:24  */
  assign n3174 = x == 10'b0000000000;
  /* fppow16.vhdl:707:24  */
  assign n3177 = x == 10'b0000000001;
  /* fppow16.vhdl:708:24  */
  assign n3180 = x == 10'b0000000010;
  /* fppow16.vhdl:709:24  */
  assign n3183 = x == 10'b0000000011;
  /* fppow16.vhdl:710:24  */
  assign n3186 = x == 10'b0000000100;
  /* fppow16.vhdl:711:24  */
  assign n3189 = x == 10'b0000000101;
  /* fppow16.vhdl:712:24  */
  assign n3192 = x == 10'b0000000110;
  /* fppow16.vhdl:713:24  */
  assign n3195 = x == 10'b0000000111;
  /* fppow16.vhdl:714:24  */
  assign n3198 = x == 10'b0000001000;
  /* fppow16.vhdl:715:24  */
  assign n3201 = x == 10'b0000001001;
  /* fppow16.vhdl:716:24  */
  assign n3204 = x == 10'b0000001010;
  /* fppow16.vhdl:717:24  */
  assign n3207 = x == 10'b0000001011;
  /* fppow16.vhdl:718:24  */
  assign n3210 = x == 10'b0000001100;
  /* fppow16.vhdl:719:24  */
  assign n3213 = x == 10'b0000001101;
  /* fppow16.vhdl:720:24  */
  assign n3216 = x == 10'b0000001110;
  /* fppow16.vhdl:721:24  */
  assign n3219 = x == 10'b0000001111;
  /* fppow16.vhdl:722:24  */
  assign n3222 = x == 10'b0000010000;
  /* fppow16.vhdl:723:24  */
  assign n3225 = x == 10'b0000010001;
  /* fppow16.vhdl:724:24  */
  assign n3228 = x == 10'b0000010010;
  /* fppow16.vhdl:725:24  */
  assign n3231 = x == 10'b0000010011;
  /* fppow16.vhdl:726:24  */
  assign n3234 = x == 10'b0000010100;
  /* fppow16.vhdl:727:24  */
  assign n3237 = x == 10'b0000010101;
  /* fppow16.vhdl:728:24  */
  assign n3240 = x == 10'b0000010110;
  /* fppow16.vhdl:729:24  */
  assign n3243 = x == 10'b0000010111;
  /* fppow16.vhdl:730:24  */
  assign n3246 = x == 10'b0000011000;
  /* fppow16.vhdl:731:24  */
  assign n3249 = x == 10'b0000011001;
  /* fppow16.vhdl:732:24  */
  assign n3252 = x == 10'b0000011010;
  /* fppow16.vhdl:733:24  */
  assign n3255 = x == 10'b0000011011;
  /* fppow16.vhdl:734:24  */
  assign n3258 = x == 10'b0000011100;
  /* fppow16.vhdl:735:24  */
  assign n3261 = x == 10'b0000011101;
  /* fppow16.vhdl:736:24  */
  assign n3264 = x == 10'b0000011110;
  /* fppow16.vhdl:737:24  */
  assign n3267 = x == 10'b0000011111;
  /* fppow16.vhdl:738:24  */
  assign n3270 = x == 10'b0000100000;
  /* fppow16.vhdl:739:24  */
  assign n3273 = x == 10'b0000100001;
  /* fppow16.vhdl:740:24  */
  assign n3276 = x == 10'b0000100010;
  /* fppow16.vhdl:741:24  */
  assign n3279 = x == 10'b0000100011;
  /* fppow16.vhdl:742:24  */
  assign n3282 = x == 10'b0000100100;
  /* fppow16.vhdl:743:24  */
  assign n3285 = x == 10'b0000100101;
  /* fppow16.vhdl:744:24  */
  assign n3288 = x == 10'b0000100110;
  /* fppow16.vhdl:745:24  */
  assign n3291 = x == 10'b0000100111;
  /* fppow16.vhdl:746:24  */
  assign n3294 = x == 10'b0000101000;
  /* fppow16.vhdl:747:24  */
  assign n3297 = x == 10'b0000101001;
  /* fppow16.vhdl:748:24  */
  assign n3300 = x == 10'b0000101010;
  /* fppow16.vhdl:749:24  */
  assign n3303 = x == 10'b0000101011;
  /* fppow16.vhdl:750:24  */
  assign n3306 = x == 10'b0000101100;
  /* fppow16.vhdl:751:24  */
  assign n3309 = x == 10'b0000101101;
  /* fppow16.vhdl:752:24  */
  assign n3312 = x == 10'b0000101110;
  /* fppow16.vhdl:753:24  */
  assign n3315 = x == 10'b0000101111;
  /* fppow16.vhdl:754:24  */
  assign n3318 = x == 10'b0000110000;
  /* fppow16.vhdl:755:24  */
  assign n3321 = x == 10'b0000110001;
  /* fppow16.vhdl:756:24  */
  assign n3324 = x == 10'b0000110010;
  /* fppow16.vhdl:757:24  */
  assign n3327 = x == 10'b0000110011;
  /* fppow16.vhdl:758:24  */
  assign n3330 = x == 10'b0000110100;
  /* fppow16.vhdl:759:24  */
  assign n3333 = x == 10'b0000110101;
  /* fppow16.vhdl:760:24  */
  assign n3336 = x == 10'b0000110110;
  /* fppow16.vhdl:761:24  */
  assign n3339 = x == 10'b0000110111;
  /* fppow16.vhdl:762:24  */
  assign n3342 = x == 10'b0000111000;
  /* fppow16.vhdl:763:24  */
  assign n3345 = x == 10'b0000111001;
  /* fppow16.vhdl:764:24  */
  assign n3348 = x == 10'b0000111010;
  /* fppow16.vhdl:765:24  */
  assign n3351 = x == 10'b0000111011;
  /* fppow16.vhdl:766:24  */
  assign n3354 = x == 10'b0000111100;
  /* fppow16.vhdl:767:24  */
  assign n3357 = x == 10'b0000111101;
  /* fppow16.vhdl:768:24  */
  assign n3360 = x == 10'b0000111110;
  /* fppow16.vhdl:769:24  */
  assign n3363 = x == 10'b0000111111;
  /* fppow16.vhdl:770:24  */
  assign n3366 = x == 10'b0001000000;
  /* fppow16.vhdl:771:24  */
  assign n3369 = x == 10'b0001000001;
  /* fppow16.vhdl:772:24  */
  assign n3372 = x == 10'b0001000010;
  /* fppow16.vhdl:773:24  */
  assign n3375 = x == 10'b0001000011;
  /* fppow16.vhdl:774:24  */
  assign n3378 = x == 10'b0001000100;
  /* fppow16.vhdl:775:24  */
  assign n3381 = x == 10'b0001000101;
  /* fppow16.vhdl:776:24  */
  assign n3384 = x == 10'b0001000110;
  /* fppow16.vhdl:777:24  */
  assign n3387 = x == 10'b0001000111;
  /* fppow16.vhdl:778:24  */
  assign n3390 = x == 10'b0001001000;
  /* fppow16.vhdl:779:24  */
  assign n3393 = x == 10'b0001001001;
  /* fppow16.vhdl:780:24  */
  assign n3396 = x == 10'b0001001010;
  /* fppow16.vhdl:781:24  */
  assign n3399 = x == 10'b0001001011;
  /* fppow16.vhdl:782:24  */
  assign n3402 = x == 10'b0001001100;
  /* fppow16.vhdl:783:24  */
  assign n3405 = x == 10'b0001001101;
  /* fppow16.vhdl:784:24  */
  assign n3408 = x == 10'b0001001110;
  /* fppow16.vhdl:785:24  */
  assign n3411 = x == 10'b0001001111;
  /* fppow16.vhdl:786:24  */
  assign n3414 = x == 10'b0001010000;
  /* fppow16.vhdl:787:24  */
  assign n3417 = x == 10'b0001010001;
  /* fppow16.vhdl:788:24  */
  assign n3420 = x == 10'b0001010010;
  /* fppow16.vhdl:789:24  */
  assign n3423 = x == 10'b0001010011;
  /* fppow16.vhdl:790:24  */
  assign n3426 = x == 10'b0001010100;
  /* fppow16.vhdl:791:24  */
  assign n3429 = x == 10'b0001010101;
  /* fppow16.vhdl:792:24  */
  assign n3432 = x == 10'b0001010110;
  /* fppow16.vhdl:793:24  */
  assign n3435 = x == 10'b0001010111;
  /* fppow16.vhdl:794:24  */
  assign n3438 = x == 10'b0001011000;
  /* fppow16.vhdl:795:24  */
  assign n3441 = x == 10'b0001011001;
  /* fppow16.vhdl:796:24  */
  assign n3444 = x == 10'b0001011010;
  /* fppow16.vhdl:797:24  */
  assign n3447 = x == 10'b0001011011;
  /* fppow16.vhdl:798:24  */
  assign n3450 = x == 10'b0001011100;
  /* fppow16.vhdl:799:24  */
  assign n3453 = x == 10'b0001011101;
  /* fppow16.vhdl:800:24  */
  assign n3456 = x == 10'b0001011110;
  /* fppow16.vhdl:801:24  */
  assign n3459 = x == 10'b0001011111;
  /* fppow16.vhdl:802:24  */
  assign n3462 = x == 10'b0001100000;
  /* fppow16.vhdl:803:24  */
  assign n3465 = x == 10'b0001100001;
  /* fppow16.vhdl:804:24  */
  assign n3468 = x == 10'b0001100010;
  /* fppow16.vhdl:805:24  */
  assign n3471 = x == 10'b0001100011;
  /* fppow16.vhdl:806:24  */
  assign n3474 = x == 10'b0001100100;
  /* fppow16.vhdl:807:24  */
  assign n3477 = x == 10'b0001100101;
  /* fppow16.vhdl:808:24  */
  assign n3480 = x == 10'b0001100110;
  /* fppow16.vhdl:809:24  */
  assign n3483 = x == 10'b0001100111;
  /* fppow16.vhdl:810:24  */
  assign n3486 = x == 10'b0001101000;
  /* fppow16.vhdl:811:24  */
  assign n3489 = x == 10'b0001101001;
  /* fppow16.vhdl:812:24  */
  assign n3492 = x == 10'b0001101010;
  /* fppow16.vhdl:813:24  */
  assign n3495 = x == 10'b0001101011;
  /* fppow16.vhdl:814:24  */
  assign n3498 = x == 10'b0001101100;
  /* fppow16.vhdl:815:24  */
  assign n3501 = x == 10'b0001101101;
  /* fppow16.vhdl:816:24  */
  assign n3504 = x == 10'b0001101110;
  /* fppow16.vhdl:817:24  */
  assign n3507 = x == 10'b0001101111;
  /* fppow16.vhdl:818:24  */
  assign n3510 = x == 10'b0001110000;
  /* fppow16.vhdl:819:24  */
  assign n3513 = x == 10'b0001110001;
  /* fppow16.vhdl:820:24  */
  assign n3516 = x == 10'b0001110010;
  /* fppow16.vhdl:821:24  */
  assign n3519 = x == 10'b0001110011;
  /* fppow16.vhdl:822:24  */
  assign n3522 = x == 10'b0001110100;
  /* fppow16.vhdl:823:24  */
  assign n3525 = x == 10'b0001110101;
  /* fppow16.vhdl:824:24  */
  assign n3528 = x == 10'b0001110110;
  /* fppow16.vhdl:825:24  */
  assign n3531 = x == 10'b0001110111;
  /* fppow16.vhdl:826:24  */
  assign n3534 = x == 10'b0001111000;
  /* fppow16.vhdl:827:24  */
  assign n3537 = x == 10'b0001111001;
  /* fppow16.vhdl:828:24  */
  assign n3540 = x == 10'b0001111010;
  /* fppow16.vhdl:829:24  */
  assign n3543 = x == 10'b0001111011;
  /* fppow16.vhdl:830:24  */
  assign n3546 = x == 10'b0001111100;
  /* fppow16.vhdl:831:24  */
  assign n3549 = x == 10'b0001111101;
  /* fppow16.vhdl:832:24  */
  assign n3552 = x == 10'b0001111110;
  /* fppow16.vhdl:833:24  */
  assign n3555 = x == 10'b0001111111;
  /* fppow16.vhdl:834:24  */
  assign n3558 = x == 10'b0010000000;
  /* fppow16.vhdl:835:24  */
  assign n3561 = x == 10'b0010000001;
  /* fppow16.vhdl:836:24  */
  assign n3564 = x == 10'b0010000010;
  /* fppow16.vhdl:837:24  */
  assign n3567 = x == 10'b0010000011;
  /* fppow16.vhdl:838:24  */
  assign n3570 = x == 10'b0010000100;
  /* fppow16.vhdl:839:24  */
  assign n3573 = x == 10'b0010000101;
  /* fppow16.vhdl:840:24  */
  assign n3576 = x == 10'b0010000110;
  /* fppow16.vhdl:841:24  */
  assign n3579 = x == 10'b0010000111;
  /* fppow16.vhdl:842:24  */
  assign n3582 = x == 10'b0010001000;
  /* fppow16.vhdl:843:24  */
  assign n3585 = x == 10'b0010001001;
  /* fppow16.vhdl:844:24  */
  assign n3588 = x == 10'b0010001010;
  /* fppow16.vhdl:845:24  */
  assign n3591 = x == 10'b0010001011;
  /* fppow16.vhdl:846:24  */
  assign n3594 = x == 10'b0010001100;
  /* fppow16.vhdl:847:24  */
  assign n3597 = x == 10'b0010001101;
  /* fppow16.vhdl:848:24  */
  assign n3600 = x == 10'b0010001110;
  /* fppow16.vhdl:849:24  */
  assign n3603 = x == 10'b0010001111;
  /* fppow16.vhdl:850:24  */
  assign n3606 = x == 10'b0010010000;
  /* fppow16.vhdl:851:24  */
  assign n3609 = x == 10'b0010010001;
  /* fppow16.vhdl:852:24  */
  assign n3612 = x == 10'b0010010010;
  /* fppow16.vhdl:853:24  */
  assign n3615 = x == 10'b0010010011;
  /* fppow16.vhdl:854:24  */
  assign n3618 = x == 10'b0010010100;
  /* fppow16.vhdl:855:24  */
  assign n3621 = x == 10'b0010010101;
  /* fppow16.vhdl:856:24  */
  assign n3624 = x == 10'b0010010110;
  /* fppow16.vhdl:857:24  */
  assign n3627 = x == 10'b0010010111;
  /* fppow16.vhdl:858:24  */
  assign n3630 = x == 10'b0010011000;
  /* fppow16.vhdl:859:24  */
  assign n3633 = x == 10'b0010011001;
  /* fppow16.vhdl:860:24  */
  assign n3636 = x == 10'b0010011010;
  /* fppow16.vhdl:861:24  */
  assign n3639 = x == 10'b0010011011;
  /* fppow16.vhdl:862:24  */
  assign n3642 = x == 10'b0010011100;
  /* fppow16.vhdl:863:24  */
  assign n3645 = x == 10'b0010011101;
  /* fppow16.vhdl:864:24  */
  assign n3648 = x == 10'b0010011110;
  /* fppow16.vhdl:865:24  */
  assign n3651 = x == 10'b0010011111;
  /* fppow16.vhdl:866:24  */
  assign n3654 = x == 10'b0010100000;
  /* fppow16.vhdl:867:24  */
  assign n3657 = x == 10'b0010100001;
  /* fppow16.vhdl:868:24  */
  assign n3660 = x == 10'b0010100010;
  /* fppow16.vhdl:869:24  */
  assign n3663 = x == 10'b0010100011;
  /* fppow16.vhdl:870:24  */
  assign n3666 = x == 10'b0010100100;
  /* fppow16.vhdl:871:24  */
  assign n3669 = x == 10'b0010100101;
  /* fppow16.vhdl:872:24  */
  assign n3672 = x == 10'b0010100110;
  /* fppow16.vhdl:873:24  */
  assign n3675 = x == 10'b0010100111;
  /* fppow16.vhdl:874:24  */
  assign n3678 = x == 10'b0010101000;
  /* fppow16.vhdl:875:24  */
  assign n3681 = x == 10'b0010101001;
  /* fppow16.vhdl:876:24  */
  assign n3684 = x == 10'b0010101010;
  /* fppow16.vhdl:877:24  */
  assign n3687 = x == 10'b0010101011;
  /* fppow16.vhdl:878:24  */
  assign n3690 = x == 10'b0010101100;
  /* fppow16.vhdl:879:24  */
  assign n3693 = x == 10'b0010101101;
  /* fppow16.vhdl:880:24  */
  assign n3696 = x == 10'b0010101110;
  /* fppow16.vhdl:881:24  */
  assign n3699 = x == 10'b0010101111;
  /* fppow16.vhdl:882:24  */
  assign n3702 = x == 10'b0010110000;
  /* fppow16.vhdl:883:24  */
  assign n3705 = x == 10'b0010110001;
  /* fppow16.vhdl:884:24  */
  assign n3708 = x == 10'b0010110010;
  /* fppow16.vhdl:885:24  */
  assign n3711 = x == 10'b0010110011;
  /* fppow16.vhdl:886:24  */
  assign n3714 = x == 10'b0010110100;
  /* fppow16.vhdl:887:24  */
  assign n3717 = x == 10'b0010110101;
  /* fppow16.vhdl:888:24  */
  assign n3720 = x == 10'b0010110110;
  /* fppow16.vhdl:889:24  */
  assign n3723 = x == 10'b0010110111;
  /* fppow16.vhdl:890:24  */
  assign n3726 = x == 10'b0010111000;
  /* fppow16.vhdl:891:24  */
  assign n3729 = x == 10'b0010111001;
  /* fppow16.vhdl:892:24  */
  assign n3732 = x == 10'b0010111010;
  /* fppow16.vhdl:893:24  */
  assign n3735 = x == 10'b0010111011;
  /* fppow16.vhdl:894:24  */
  assign n3738 = x == 10'b0010111100;
  /* fppow16.vhdl:895:24  */
  assign n3741 = x == 10'b0010111101;
  /* fppow16.vhdl:896:24  */
  assign n3744 = x == 10'b0010111110;
  /* fppow16.vhdl:897:24  */
  assign n3747 = x == 10'b0010111111;
  /* fppow16.vhdl:898:24  */
  assign n3750 = x == 10'b0011000000;
  /* fppow16.vhdl:899:24  */
  assign n3753 = x == 10'b0011000001;
  /* fppow16.vhdl:900:24  */
  assign n3756 = x == 10'b0011000010;
  /* fppow16.vhdl:901:24  */
  assign n3759 = x == 10'b0011000011;
  /* fppow16.vhdl:902:24  */
  assign n3762 = x == 10'b0011000100;
  /* fppow16.vhdl:903:24  */
  assign n3765 = x == 10'b0011000101;
  /* fppow16.vhdl:904:24  */
  assign n3768 = x == 10'b0011000110;
  /* fppow16.vhdl:905:24  */
  assign n3771 = x == 10'b0011000111;
  /* fppow16.vhdl:906:24  */
  assign n3774 = x == 10'b0011001000;
  /* fppow16.vhdl:907:24  */
  assign n3777 = x == 10'b0011001001;
  /* fppow16.vhdl:908:24  */
  assign n3780 = x == 10'b0011001010;
  /* fppow16.vhdl:909:24  */
  assign n3783 = x == 10'b0011001011;
  /* fppow16.vhdl:910:24  */
  assign n3786 = x == 10'b0011001100;
  /* fppow16.vhdl:911:24  */
  assign n3789 = x == 10'b0011001101;
  /* fppow16.vhdl:912:24  */
  assign n3792 = x == 10'b0011001110;
  /* fppow16.vhdl:913:24  */
  assign n3795 = x == 10'b0011001111;
  /* fppow16.vhdl:914:24  */
  assign n3798 = x == 10'b0011010000;
  /* fppow16.vhdl:915:24  */
  assign n3801 = x == 10'b0011010001;
  /* fppow16.vhdl:916:24  */
  assign n3804 = x == 10'b0011010010;
  /* fppow16.vhdl:917:24  */
  assign n3807 = x == 10'b0011010011;
  /* fppow16.vhdl:918:24  */
  assign n3810 = x == 10'b0011010100;
  /* fppow16.vhdl:919:24  */
  assign n3813 = x == 10'b0011010101;
  /* fppow16.vhdl:920:24  */
  assign n3816 = x == 10'b0011010110;
  /* fppow16.vhdl:921:24  */
  assign n3819 = x == 10'b0011010111;
  /* fppow16.vhdl:922:24  */
  assign n3822 = x == 10'b0011011000;
  /* fppow16.vhdl:923:24  */
  assign n3825 = x == 10'b0011011001;
  /* fppow16.vhdl:924:24  */
  assign n3828 = x == 10'b0011011010;
  /* fppow16.vhdl:925:24  */
  assign n3831 = x == 10'b0011011011;
  /* fppow16.vhdl:926:24  */
  assign n3834 = x == 10'b0011011100;
  /* fppow16.vhdl:927:24  */
  assign n3837 = x == 10'b0011011101;
  /* fppow16.vhdl:928:24  */
  assign n3840 = x == 10'b0011011110;
  /* fppow16.vhdl:929:24  */
  assign n3843 = x == 10'b0011011111;
  /* fppow16.vhdl:930:24  */
  assign n3846 = x == 10'b0011100000;
  /* fppow16.vhdl:931:24  */
  assign n3849 = x == 10'b0011100001;
  /* fppow16.vhdl:932:24  */
  assign n3852 = x == 10'b0011100010;
  /* fppow16.vhdl:933:24  */
  assign n3855 = x == 10'b0011100011;
  /* fppow16.vhdl:934:24  */
  assign n3858 = x == 10'b0011100100;
  /* fppow16.vhdl:935:24  */
  assign n3861 = x == 10'b0011100101;
  /* fppow16.vhdl:936:24  */
  assign n3864 = x == 10'b0011100110;
  /* fppow16.vhdl:937:24  */
  assign n3867 = x == 10'b0011100111;
  /* fppow16.vhdl:938:24  */
  assign n3870 = x == 10'b0011101000;
  /* fppow16.vhdl:939:24  */
  assign n3873 = x == 10'b0011101001;
  /* fppow16.vhdl:940:24  */
  assign n3876 = x == 10'b0011101010;
  /* fppow16.vhdl:941:24  */
  assign n3879 = x == 10'b0011101011;
  /* fppow16.vhdl:942:24  */
  assign n3882 = x == 10'b0011101100;
  /* fppow16.vhdl:943:24  */
  assign n3885 = x == 10'b0011101101;
  /* fppow16.vhdl:944:24  */
  assign n3888 = x == 10'b0011101110;
  /* fppow16.vhdl:945:24  */
  assign n3891 = x == 10'b0011101111;
  /* fppow16.vhdl:946:24  */
  assign n3894 = x == 10'b0011110000;
  /* fppow16.vhdl:947:24  */
  assign n3897 = x == 10'b0011110001;
  /* fppow16.vhdl:948:24  */
  assign n3900 = x == 10'b0011110010;
  /* fppow16.vhdl:949:24  */
  assign n3903 = x == 10'b0011110011;
  /* fppow16.vhdl:950:24  */
  assign n3906 = x == 10'b0011110100;
  /* fppow16.vhdl:951:24  */
  assign n3909 = x == 10'b0011110101;
  /* fppow16.vhdl:952:24  */
  assign n3912 = x == 10'b0011110110;
  /* fppow16.vhdl:953:24  */
  assign n3915 = x == 10'b0011110111;
  /* fppow16.vhdl:954:24  */
  assign n3918 = x == 10'b0011111000;
  /* fppow16.vhdl:955:24  */
  assign n3921 = x == 10'b0011111001;
  /* fppow16.vhdl:956:24  */
  assign n3924 = x == 10'b0011111010;
  /* fppow16.vhdl:957:24  */
  assign n3927 = x == 10'b0011111011;
  /* fppow16.vhdl:958:24  */
  assign n3930 = x == 10'b0011111100;
  /* fppow16.vhdl:959:24  */
  assign n3933 = x == 10'b0011111101;
  /* fppow16.vhdl:960:24  */
  assign n3936 = x == 10'b0011111110;
  /* fppow16.vhdl:961:24  */
  assign n3939 = x == 10'b0011111111;
  /* fppow16.vhdl:962:24  */
  assign n3942 = x == 10'b0100000000;
  /* fppow16.vhdl:963:24  */
  assign n3945 = x == 10'b0100000001;
  /* fppow16.vhdl:964:24  */
  assign n3948 = x == 10'b0100000010;
  /* fppow16.vhdl:965:24  */
  assign n3951 = x == 10'b0100000011;
  /* fppow16.vhdl:966:24  */
  assign n3954 = x == 10'b0100000100;
  /* fppow16.vhdl:967:24  */
  assign n3957 = x == 10'b0100000101;
  /* fppow16.vhdl:968:24  */
  assign n3960 = x == 10'b0100000110;
  /* fppow16.vhdl:969:24  */
  assign n3963 = x == 10'b0100000111;
  /* fppow16.vhdl:970:24  */
  assign n3966 = x == 10'b0100001000;
  /* fppow16.vhdl:971:24  */
  assign n3969 = x == 10'b0100001001;
  /* fppow16.vhdl:972:24  */
  assign n3972 = x == 10'b0100001010;
  /* fppow16.vhdl:973:24  */
  assign n3975 = x == 10'b0100001011;
  /* fppow16.vhdl:974:24  */
  assign n3978 = x == 10'b0100001100;
  /* fppow16.vhdl:975:24  */
  assign n3981 = x == 10'b0100001101;
  /* fppow16.vhdl:976:24  */
  assign n3984 = x == 10'b0100001110;
  /* fppow16.vhdl:977:24  */
  assign n3987 = x == 10'b0100001111;
  /* fppow16.vhdl:978:24  */
  assign n3990 = x == 10'b0100010000;
  /* fppow16.vhdl:979:24  */
  assign n3993 = x == 10'b0100010001;
  /* fppow16.vhdl:980:24  */
  assign n3996 = x == 10'b0100010010;
  /* fppow16.vhdl:981:24  */
  assign n3999 = x == 10'b0100010011;
  /* fppow16.vhdl:982:24  */
  assign n4002 = x == 10'b0100010100;
  /* fppow16.vhdl:983:24  */
  assign n4005 = x == 10'b0100010101;
  /* fppow16.vhdl:984:24  */
  assign n4008 = x == 10'b0100010110;
  /* fppow16.vhdl:985:24  */
  assign n4011 = x == 10'b0100010111;
  /* fppow16.vhdl:986:24  */
  assign n4014 = x == 10'b0100011000;
  /* fppow16.vhdl:987:24  */
  assign n4017 = x == 10'b0100011001;
  /* fppow16.vhdl:988:24  */
  assign n4020 = x == 10'b0100011010;
  /* fppow16.vhdl:989:24  */
  assign n4023 = x == 10'b0100011011;
  /* fppow16.vhdl:990:24  */
  assign n4026 = x == 10'b0100011100;
  /* fppow16.vhdl:991:24  */
  assign n4029 = x == 10'b0100011101;
  /* fppow16.vhdl:992:24  */
  assign n4032 = x == 10'b0100011110;
  /* fppow16.vhdl:993:24  */
  assign n4035 = x == 10'b0100011111;
  /* fppow16.vhdl:994:24  */
  assign n4038 = x == 10'b0100100000;
  /* fppow16.vhdl:995:24  */
  assign n4041 = x == 10'b0100100001;
  /* fppow16.vhdl:996:24  */
  assign n4044 = x == 10'b0100100010;
  /* fppow16.vhdl:997:24  */
  assign n4047 = x == 10'b0100100011;
  /* fppow16.vhdl:998:24  */
  assign n4050 = x == 10'b0100100100;
  /* fppow16.vhdl:999:24  */
  assign n4053 = x == 10'b0100100101;
  /* fppow16.vhdl:1000:24  */
  assign n4056 = x == 10'b0100100110;
  /* fppow16.vhdl:1001:24  */
  assign n4059 = x == 10'b0100100111;
  /* fppow16.vhdl:1002:24  */
  assign n4062 = x == 10'b0100101000;
  /* fppow16.vhdl:1003:24  */
  assign n4065 = x == 10'b0100101001;
  /* fppow16.vhdl:1004:24  */
  assign n4068 = x == 10'b0100101010;
  /* fppow16.vhdl:1005:24  */
  assign n4071 = x == 10'b0100101011;
  /* fppow16.vhdl:1006:24  */
  assign n4074 = x == 10'b0100101100;
  /* fppow16.vhdl:1007:24  */
  assign n4077 = x == 10'b0100101101;
  /* fppow16.vhdl:1008:24  */
  assign n4080 = x == 10'b0100101110;
  /* fppow16.vhdl:1009:24  */
  assign n4083 = x == 10'b0100101111;
  /* fppow16.vhdl:1010:24  */
  assign n4086 = x == 10'b0100110000;
  /* fppow16.vhdl:1011:24  */
  assign n4089 = x == 10'b0100110001;
  /* fppow16.vhdl:1012:24  */
  assign n4092 = x == 10'b0100110010;
  /* fppow16.vhdl:1013:24  */
  assign n4095 = x == 10'b0100110011;
  /* fppow16.vhdl:1014:24  */
  assign n4098 = x == 10'b0100110100;
  /* fppow16.vhdl:1015:24  */
  assign n4101 = x == 10'b0100110101;
  /* fppow16.vhdl:1016:24  */
  assign n4104 = x == 10'b0100110110;
  /* fppow16.vhdl:1017:24  */
  assign n4107 = x == 10'b0100110111;
  /* fppow16.vhdl:1018:24  */
  assign n4110 = x == 10'b0100111000;
  /* fppow16.vhdl:1019:24  */
  assign n4113 = x == 10'b0100111001;
  /* fppow16.vhdl:1020:24  */
  assign n4116 = x == 10'b0100111010;
  /* fppow16.vhdl:1021:24  */
  assign n4119 = x == 10'b0100111011;
  /* fppow16.vhdl:1022:24  */
  assign n4122 = x == 10'b0100111100;
  /* fppow16.vhdl:1023:24  */
  assign n4125 = x == 10'b0100111101;
  /* fppow16.vhdl:1024:24  */
  assign n4128 = x == 10'b0100111110;
  /* fppow16.vhdl:1025:24  */
  assign n4131 = x == 10'b0100111111;
  /* fppow16.vhdl:1026:24  */
  assign n4134 = x == 10'b0101000000;
  /* fppow16.vhdl:1027:24  */
  assign n4137 = x == 10'b0101000001;
  /* fppow16.vhdl:1028:24  */
  assign n4140 = x == 10'b0101000010;
  /* fppow16.vhdl:1029:24  */
  assign n4143 = x == 10'b0101000011;
  /* fppow16.vhdl:1030:24  */
  assign n4146 = x == 10'b0101000100;
  /* fppow16.vhdl:1031:24  */
  assign n4149 = x == 10'b0101000101;
  /* fppow16.vhdl:1032:24  */
  assign n4152 = x == 10'b0101000110;
  /* fppow16.vhdl:1033:24  */
  assign n4155 = x == 10'b0101000111;
  /* fppow16.vhdl:1034:24  */
  assign n4158 = x == 10'b0101001000;
  /* fppow16.vhdl:1035:24  */
  assign n4161 = x == 10'b0101001001;
  /* fppow16.vhdl:1036:24  */
  assign n4164 = x == 10'b0101001010;
  /* fppow16.vhdl:1037:24  */
  assign n4167 = x == 10'b0101001011;
  /* fppow16.vhdl:1038:24  */
  assign n4170 = x == 10'b0101001100;
  /* fppow16.vhdl:1039:24  */
  assign n4173 = x == 10'b0101001101;
  /* fppow16.vhdl:1040:24  */
  assign n4176 = x == 10'b0101001110;
  /* fppow16.vhdl:1041:24  */
  assign n4179 = x == 10'b0101001111;
  /* fppow16.vhdl:1042:24  */
  assign n4182 = x == 10'b0101010000;
  /* fppow16.vhdl:1043:24  */
  assign n4185 = x == 10'b0101010001;
  /* fppow16.vhdl:1044:24  */
  assign n4188 = x == 10'b0101010010;
  /* fppow16.vhdl:1045:24  */
  assign n4191 = x == 10'b0101010011;
  /* fppow16.vhdl:1046:24  */
  assign n4194 = x == 10'b0101010100;
  /* fppow16.vhdl:1047:24  */
  assign n4197 = x == 10'b0101010101;
  /* fppow16.vhdl:1048:24  */
  assign n4200 = x == 10'b0101010110;
  /* fppow16.vhdl:1049:24  */
  assign n4203 = x == 10'b0101010111;
  /* fppow16.vhdl:1050:24  */
  assign n4206 = x == 10'b0101011000;
  /* fppow16.vhdl:1051:24  */
  assign n4209 = x == 10'b0101011001;
  /* fppow16.vhdl:1052:24  */
  assign n4212 = x == 10'b0101011010;
  /* fppow16.vhdl:1053:24  */
  assign n4215 = x == 10'b0101011011;
  /* fppow16.vhdl:1054:24  */
  assign n4218 = x == 10'b0101011100;
  /* fppow16.vhdl:1055:24  */
  assign n4221 = x == 10'b0101011101;
  /* fppow16.vhdl:1056:24  */
  assign n4224 = x == 10'b0101011110;
  /* fppow16.vhdl:1057:24  */
  assign n4227 = x == 10'b0101011111;
  /* fppow16.vhdl:1058:24  */
  assign n4230 = x == 10'b0101100000;
  /* fppow16.vhdl:1059:24  */
  assign n4233 = x == 10'b0101100001;
  /* fppow16.vhdl:1060:24  */
  assign n4236 = x == 10'b0101100010;
  /* fppow16.vhdl:1061:24  */
  assign n4239 = x == 10'b0101100011;
  /* fppow16.vhdl:1062:24  */
  assign n4242 = x == 10'b0101100100;
  /* fppow16.vhdl:1063:24  */
  assign n4245 = x == 10'b0101100101;
  /* fppow16.vhdl:1064:24  */
  assign n4248 = x == 10'b0101100110;
  /* fppow16.vhdl:1065:24  */
  assign n4251 = x == 10'b0101100111;
  /* fppow16.vhdl:1066:24  */
  assign n4254 = x == 10'b0101101000;
  /* fppow16.vhdl:1067:24  */
  assign n4257 = x == 10'b0101101001;
  /* fppow16.vhdl:1068:24  */
  assign n4260 = x == 10'b0101101010;
  /* fppow16.vhdl:1069:24  */
  assign n4263 = x == 10'b0101101011;
  /* fppow16.vhdl:1070:24  */
  assign n4266 = x == 10'b0101101100;
  /* fppow16.vhdl:1071:24  */
  assign n4269 = x == 10'b0101101101;
  /* fppow16.vhdl:1072:24  */
  assign n4272 = x == 10'b0101101110;
  /* fppow16.vhdl:1073:24  */
  assign n4275 = x == 10'b0101101111;
  /* fppow16.vhdl:1074:24  */
  assign n4278 = x == 10'b0101110000;
  /* fppow16.vhdl:1075:24  */
  assign n4281 = x == 10'b0101110001;
  /* fppow16.vhdl:1076:24  */
  assign n4284 = x == 10'b0101110010;
  /* fppow16.vhdl:1077:24  */
  assign n4287 = x == 10'b0101110011;
  /* fppow16.vhdl:1078:24  */
  assign n4290 = x == 10'b0101110100;
  /* fppow16.vhdl:1079:24  */
  assign n4293 = x == 10'b0101110101;
  /* fppow16.vhdl:1080:24  */
  assign n4296 = x == 10'b0101110110;
  /* fppow16.vhdl:1081:24  */
  assign n4299 = x == 10'b0101110111;
  /* fppow16.vhdl:1082:24  */
  assign n4302 = x == 10'b0101111000;
  /* fppow16.vhdl:1083:24  */
  assign n4305 = x == 10'b0101111001;
  /* fppow16.vhdl:1084:24  */
  assign n4308 = x == 10'b0101111010;
  /* fppow16.vhdl:1085:24  */
  assign n4311 = x == 10'b0101111011;
  /* fppow16.vhdl:1086:24  */
  assign n4314 = x == 10'b0101111100;
  /* fppow16.vhdl:1087:24  */
  assign n4317 = x == 10'b0101111101;
  /* fppow16.vhdl:1088:24  */
  assign n4320 = x == 10'b0101111110;
  /* fppow16.vhdl:1089:24  */
  assign n4323 = x == 10'b0101111111;
  /* fppow16.vhdl:1090:24  */
  assign n4326 = x == 10'b0110000000;
  /* fppow16.vhdl:1091:24  */
  assign n4329 = x == 10'b0110000001;
  /* fppow16.vhdl:1092:24  */
  assign n4332 = x == 10'b0110000010;
  /* fppow16.vhdl:1093:24  */
  assign n4335 = x == 10'b0110000011;
  /* fppow16.vhdl:1094:24  */
  assign n4338 = x == 10'b0110000100;
  /* fppow16.vhdl:1095:24  */
  assign n4341 = x == 10'b0110000101;
  /* fppow16.vhdl:1096:24  */
  assign n4344 = x == 10'b0110000110;
  /* fppow16.vhdl:1097:24  */
  assign n4347 = x == 10'b0110000111;
  /* fppow16.vhdl:1098:24  */
  assign n4350 = x == 10'b0110001000;
  /* fppow16.vhdl:1099:24  */
  assign n4353 = x == 10'b0110001001;
  /* fppow16.vhdl:1100:24  */
  assign n4356 = x == 10'b0110001010;
  /* fppow16.vhdl:1101:24  */
  assign n4359 = x == 10'b0110001011;
  /* fppow16.vhdl:1102:24  */
  assign n4362 = x == 10'b0110001100;
  /* fppow16.vhdl:1103:24  */
  assign n4365 = x == 10'b0110001101;
  /* fppow16.vhdl:1104:24  */
  assign n4368 = x == 10'b0110001110;
  /* fppow16.vhdl:1105:24  */
  assign n4371 = x == 10'b0110001111;
  /* fppow16.vhdl:1106:24  */
  assign n4374 = x == 10'b0110010000;
  /* fppow16.vhdl:1107:24  */
  assign n4377 = x == 10'b0110010001;
  /* fppow16.vhdl:1108:24  */
  assign n4380 = x == 10'b0110010010;
  /* fppow16.vhdl:1109:24  */
  assign n4383 = x == 10'b0110010011;
  /* fppow16.vhdl:1110:24  */
  assign n4386 = x == 10'b0110010100;
  /* fppow16.vhdl:1111:24  */
  assign n4389 = x == 10'b0110010101;
  /* fppow16.vhdl:1112:24  */
  assign n4392 = x == 10'b0110010110;
  /* fppow16.vhdl:1113:24  */
  assign n4395 = x == 10'b0110010111;
  /* fppow16.vhdl:1114:24  */
  assign n4398 = x == 10'b0110011000;
  /* fppow16.vhdl:1115:24  */
  assign n4401 = x == 10'b0110011001;
  /* fppow16.vhdl:1116:24  */
  assign n4404 = x == 10'b0110011010;
  /* fppow16.vhdl:1117:24  */
  assign n4407 = x == 10'b0110011011;
  /* fppow16.vhdl:1118:24  */
  assign n4410 = x == 10'b0110011100;
  /* fppow16.vhdl:1119:24  */
  assign n4413 = x == 10'b0110011101;
  /* fppow16.vhdl:1120:24  */
  assign n4416 = x == 10'b0110011110;
  /* fppow16.vhdl:1121:24  */
  assign n4419 = x == 10'b0110011111;
  /* fppow16.vhdl:1122:24  */
  assign n4422 = x == 10'b0110100000;
  /* fppow16.vhdl:1123:24  */
  assign n4425 = x == 10'b0110100001;
  /* fppow16.vhdl:1124:24  */
  assign n4428 = x == 10'b0110100010;
  /* fppow16.vhdl:1125:24  */
  assign n4431 = x == 10'b0110100011;
  /* fppow16.vhdl:1126:24  */
  assign n4434 = x == 10'b0110100100;
  /* fppow16.vhdl:1127:24  */
  assign n4437 = x == 10'b0110100101;
  /* fppow16.vhdl:1128:24  */
  assign n4440 = x == 10'b0110100110;
  /* fppow16.vhdl:1129:24  */
  assign n4443 = x == 10'b0110100111;
  /* fppow16.vhdl:1130:24  */
  assign n4446 = x == 10'b0110101000;
  /* fppow16.vhdl:1131:24  */
  assign n4449 = x == 10'b0110101001;
  /* fppow16.vhdl:1132:24  */
  assign n4452 = x == 10'b0110101010;
  /* fppow16.vhdl:1133:24  */
  assign n4455 = x == 10'b0110101011;
  /* fppow16.vhdl:1134:24  */
  assign n4458 = x == 10'b0110101100;
  /* fppow16.vhdl:1135:24  */
  assign n4461 = x == 10'b0110101101;
  /* fppow16.vhdl:1136:24  */
  assign n4464 = x == 10'b0110101110;
  /* fppow16.vhdl:1137:24  */
  assign n4467 = x == 10'b0110101111;
  /* fppow16.vhdl:1138:24  */
  assign n4470 = x == 10'b0110110000;
  /* fppow16.vhdl:1139:24  */
  assign n4473 = x == 10'b0110110001;
  /* fppow16.vhdl:1140:24  */
  assign n4476 = x == 10'b0110110010;
  /* fppow16.vhdl:1141:24  */
  assign n4479 = x == 10'b0110110011;
  /* fppow16.vhdl:1142:24  */
  assign n4482 = x == 10'b0110110100;
  /* fppow16.vhdl:1143:24  */
  assign n4485 = x == 10'b0110110101;
  /* fppow16.vhdl:1144:24  */
  assign n4488 = x == 10'b0110110110;
  /* fppow16.vhdl:1145:24  */
  assign n4491 = x == 10'b0110110111;
  /* fppow16.vhdl:1146:24  */
  assign n4494 = x == 10'b0110111000;
  /* fppow16.vhdl:1147:24  */
  assign n4497 = x == 10'b0110111001;
  /* fppow16.vhdl:1148:24  */
  assign n4500 = x == 10'b0110111010;
  /* fppow16.vhdl:1149:24  */
  assign n4503 = x == 10'b0110111011;
  /* fppow16.vhdl:1150:24  */
  assign n4506 = x == 10'b0110111100;
  /* fppow16.vhdl:1151:24  */
  assign n4509 = x == 10'b0110111101;
  /* fppow16.vhdl:1152:24  */
  assign n4512 = x == 10'b0110111110;
  /* fppow16.vhdl:1153:24  */
  assign n4515 = x == 10'b0110111111;
  /* fppow16.vhdl:1154:24  */
  assign n4518 = x == 10'b0111000000;
  /* fppow16.vhdl:1155:24  */
  assign n4521 = x == 10'b0111000001;
  /* fppow16.vhdl:1156:24  */
  assign n4524 = x == 10'b0111000010;
  /* fppow16.vhdl:1157:24  */
  assign n4527 = x == 10'b0111000011;
  /* fppow16.vhdl:1158:24  */
  assign n4530 = x == 10'b0111000100;
  /* fppow16.vhdl:1159:24  */
  assign n4533 = x == 10'b0111000101;
  /* fppow16.vhdl:1160:24  */
  assign n4536 = x == 10'b0111000110;
  /* fppow16.vhdl:1161:24  */
  assign n4539 = x == 10'b0111000111;
  /* fppow16.vhdl:1162:24  */
  assign n4542 = x == 10'b0111001000;
  /* fppow16.vhdl:1163:24  */
  assign n4545 = x == 10'b0111001001;
  /* fppow16.vhdl:1164:24  */
  assign n4548 = x == 10'b0111001010;
  /* fppow16.vhdl:1165:24  */
  assign n4551 = x == 10'b0111001011;
  /* fppow16.vhdl:1166:24  */
  assign n4554 = x == 10'b0111001100;
  /* fppow16.vhdl:1167:24  */
  assign n4557 = x == 10'b0111001101;
  /* fppow16.vhdl:1168:24  */
  assign n4560 = x == 10'b0111001110;
  /* fppow16.vhdl:1169:24  */
  assign n4563 = x == 10'b0111001111;
  /* fppow16.vhdl:1170:24  */
  assign n4566 = x == 10'b0111010000;
  /* fppow16.vhdl:1171:24  */
  assign n4569 = x == 10'b0111010001;
  /* fppow16.vhdl:1172:24  */
  assign n4572 = x == 10'b0111010010;
  /* fppow16.vhdl:1173:24  */
  assign n4575 = x == 10'b0111010011;
  /* fppow16.vhdl:1174:24  */
  assign n4578 = x == 10'b0111010100;
  /* fppow16.vhdl:1175:24  */
  assign n4581 = x == 10'b0111010101;
  /* fppow16.vhdl:1176:24  */
  assign n4584 = x == 10'b0111010110;
  /* fppow16.vhdl:1177:24  */
  assign n4587 = x == 10'b0111010111;
  /* fppow16.vhdl:1178:24  */
  assign n4590 = x == 10'b0111011000;
  /* fppow16.vhdl:1179:24  */
  assign n4593 = x == 10'b0111011001;
  /* fppow16.vhdl:1180:24  */
  assign n4596 = x == 10'b0111011010;
  /* fppow16.vhdl:1181:24  */
  assign n4599 = x == 10'b0111011011;
  /* fppow16.vhdl:1182:24  */
  assign n4602 = x == 10'b0111011100;
  /* fppow16.vhdl:1183:24  */
  assign n4605 = x == 10'b0111011101;
  /* fppow16.vhdl:1184:24  */
  assign n4608 = x == 10'b0111011110;
  /* fppow16.vhdl:1185:24  */
  assign n4611 = x == 10'b0111011111;
  /* fppow16.vhdl:1186:24  */
  assign n4614 = x == 10'b0111100000;
  /* fppow16.vhdl:1187:24  */
  assign n4617 = x == 10'b0111100001;
  /* fppow16.vhdl:1188:24  */
  assign n4620 = x == 10'b0111100010;
  /* fppow16.vhdl:1189:24  */
  assign n4623 = x == 10'b0111100011;
  /* fppow16.vhdl:1190:24  */
  assign n4626 = x == 10'b0111100100;
  /* fppow16.vhdl:1191:24  */
  assign n4629 = x == 10'b0111100101;
  /* fppow16.vhdl:1192:24  */
  assign n4632 = x == 10'b0111100110;
  /* fppow16.vhdl:1193:24  */
  assign n4635 = x == 10'b0111100111;
  /* fppow16.vhdl:1194:24  */
  assign n4638 = x == 10'b0111101000;
  /* fppow16.vhdl:1195:24  */
  assign n4641 = x == 10'b0111101001;
  /* fppow16.vhdl:1196:24  */
  assign n4644 = x == 10'b0111101010;
  /* fppow16.vhdl:1197:24  */
  assign n4647 = x == 10'b0111101011;
  /* fppow16.vhdl:1198:24  */
  assign n4650 = x == 10'b0111101100;
  /* fppow16.vhdl:1199:24  */
  assign n4653 = x == 10'b0111101101;
  /* fppow16.vhdl:1200:24  */
  assign n4656 = x == 10'b0111101110;
  /* fppow16.vhdl:1201:24  */
  assign n4659 = x == 10'b0111101111;
  /* fppow16.vhdl:1202:24  */
  assign n4662 = x == 10'b0111110000;
  /* fppow16.vhdl:1203:24  */
  assign n4665 = x == 10'b0111110001;
  /* fppow16.vhdl:1204:24  */
  assign n4668 = x == 10'b0111110010;
  /* fppow16.vhdl:1205:24  */
  assign n4671 = x == 10'b0111110011;
  /* fppow16.vhdl:1206:24  */
  assign n4674 = x == 10'b0111110100;
  /* fppow16.vhdl:1207:24  */
  assign n4677 = x == 10'b0111110101;
  /* fppow16.vhdl:1208:24  */
  assign n4680 = x == 10'b0111110110;
  /* fppow16.vhdl:1209:24  */
  assign n4683 = x == 10'b0111110111;
  /* fppow16.vhdl:1210:24  */
  assign n4686 = x == 10'b0111111000;
  /* fppow16.vhdl:1211:24  */
  assign n4689 = x == 10'b0111111001;
  /* fppow16.vhdl:1212:24  */
  assign n4692 = x == 10'b0111111010;
  /* fppow16.vhdl:1213:24  */
  assign n4695 = x == 10'b0111111011;
  /* fppow16.vhdl:1214:24  */
  assign n4698 = x == 10'b0111111100;
  /* fppow16.vhdl:1215:24  */
  assign n4701 = x == 10'b0111111101;
  /* fppow16.vhdl:1216:24  */
  assign n4704 = x == 10'b0111111110;
  /* fppow16.vhdl:1217:24  */
  assign n4707 = x == 10'b0111111111;
  /* fppow16.vhdl:1218:24  */
  assign n4710 = x == 10'b1000000000;
  /* fppow16.vhdl:1219:24  */
  assign n4713 = x == 10'b1000000001;
  /* fppow16.vhdl:1220:24  */
  assign n4716 = x == 10'b1000000010;
  /* fppow16.vhdl:1221:24  */
  assign n4719 = x == 10'b1000000011;
  /* fppow16.vhdl:1222:24  */
  assign n4722 = x == 10'b1000000100;
  /* fppow16.vhdl:1223:24  */
  assign n4725 = x == 10'b1000000101;
  /* fppow16.vhdl:1224:24  */
  assign n4728 = x == 10'b1000000110;
  /* fppow16.vhdl:1225:24  */
  assign n4731 = x == 10'b1000000111;
  /* fppow16.vhdl:1226:24  */
  assign n4734 = x == 10'b1000001000;
  /* fppow16.vhdl:1227:24  */
  assign n4737 = x == 10'b1000001001;
  /* fppow16.vhdl:1228:24  */
  assign n4740 = x == 10'b1000001010;
  /* fppow16.vhdl:1229:24  */
  assign n4743 = x == 10'b1000001011;
  /* fppow16.vhdl:1230:24  */
  assign n4746 = x == 10'b1000001100;
  /* fppow16.vhdl:1231:24  */
  assign n4749 = x == 10'b1000001101;
  /* fppow16.vhdl:1232:24  */
  assign n4752 = x == 10'b1000001110;
  /* fppow16.vhdl:1233:24  */
  assign n4755 = x == 10'b1000001111;
  /* fppow16.vhdl:1234:24  */
  assign n4758 = x == 10'b1000010000;
  /* fppow16.vhdl:1235:24  */
  assign n4761 = x == 10'b1000010001;
  /* fppow16.vhdl:1236:24  */
  assign n4764 = x == 10'b1000010010;
  /* fppow16.vhdl:1237:24  */
  assign n4767 = x == 10'b1000010011;
  /* fppow16.vhdl:1238:24  */
  assign n4770 = x == 10'b1000010100;
  /* fppow16.vhdl:1239:24  */
  assign n4773 = x == 10'b1000010101;
  /* fppow16.vhdl:1240:24  */
  assign n4776 = x == 10'b1000010110;
  /* fppow16.vhdl:1241:24  */
  assign n4779 = x == 10'b1000010111;
  /* fppow16.vhdl:1242:24  */
  assign n4782 = x == 10'b1000011000;
  /* fppow16.vhdl:1243:24  */
  assign n4785 = x == 10'b1000011001;
  /* fppow16.vhdl:1244:24  */
  assign n4788 = x == 10'b1000011010;
  /* fppow16.vhdl:1245:24  */
  assign n4791 = x == 10'b1000011011;
  /* fppow16.vhdl:1246:24  */
  assign n4794 = x == 10'b1000011100;
  /* fppow16.vhdl:1247:24  */
  assign n4797 = x == 10'b1000011101;
  /* fppow16.vhdl:1248:24  */
  assign n4800 = x == 10'b1000011110;
  /* fppow16.vhdl:1249:24  */
  assign n4803 = x == 10'b1000011111;
  /* fppow16.vhdl:1250:24  */
  assign n4806 = x == 10'b1000100000;
  /* fppow16.vhdl:1251:24  */
  assign n4809 = x == 10'b1000100001;
  /* fppow16.vhdl:1252:24  */
  assign n4812 = x == 10'b1000100010;
  /* fppow16.vhdl:1253:24  */
  assign n4815 = x == 10'b1000100011;
  /* fppow16.vhdl:1254:24  */
  assign n4818 = x == 10'b1000100100;
  /* fppow16.vhdl:1255:24  */
  assign n4821 = x == 10'b1000100101;
  /* fppow16.vhdl:1256:24  */
  assign n4824 = x == 10'b1000100110;
  /* fppow16.vhdl:1257:24  */
  assign n4827 = x == 10'b1000100111;
  /* fppow16.vhdl:1258:24  */
  assign n4830 = x == 10'b1000101000;
  /* fppow16.vhdl:1259:24  */
  assign n4833 = x == 10'b1000101001;
  /* fppow16.vhdl:1260:24  */
  assign n4836 = x == 10'b1000101010;
  /* fppow16.vhdl:1261:24  */
  assign n4839 = x == 10'b1000101011;
  /* fppow16.vhdl:1262:24  */
  assign n4842 = x == 10'b1000101100;
  /* fppow16.vhdl:1263:24  */
  assign n4845 = x == 10'b1000101101;
  /* fppow16.vhdl:1264:24  */
  assign n4848 = x == 10'b1000101110;
  /* fppow16.vhdl:1265:24  */
  assign n4851 = x == 10'b1000101111;
  /* fppow16.vhdl:1266:24  */
  assign n4854 = x == 10'b1000110000;
  /* fppow16.vhdl:1267:24  */
  assign n4857 = x == 10'b1000110001;
  /* fppow16.vhdl:1268:24  */
  assign n4860 = x == 10'b1000110010;
  /* fppow16.vhdl:1269:24  */
  assign n4863 = x == 10'b1000110011;
  /* fppow16.vhdl:1270:24  */
  assign n4866 = x == 10'b1000110100;
  /* fppow16.vhdl:1271:24  */
  assign n4869 = x == 10'b1000110101;
  /* fppow16.vhdl:1272:24  */
  assign n4872 = x == 10'b1000110110;
  /* fppow16.vhdl:1273:24  */
  assign n4875 = x == 10'b1000110111;
  /* fppow16.vhdl:1274:24  */
  assign n4878 = x == 10'b1000111000;
  /* fppow16.vhdl:1275:24  */
  assign n4881 = x == 10'b1000111001;
  /* fppow16.vhdl:1276:24  */
  assign n4884 = x == 10'b1000111010;
  /* fppow16.vhdl:1277:24  */
  assign n4887 = x == 10'b1000111011;
  /* fppow16.vhdl:1278:24  */
  assign n4890 = x == 10'b1000111100;
  /* fppow16.vhdl:1279:24  */
  assign n4893 = x == 10'b1000111101;
  /* fppow16.vhdl:1280:24  */
  assign n4896 = x == 10'b1000111110;
  /* fppow16.vhdl:1281:24  */
  assign n4899 = x == 10'b1000111111;
  /* fppow16.vhdl:1282:24  */
  assign n4902 = x == 10'b1001000000;
  /* fppow16.vhdl:1283:24  */
  assign n4905 = x == 10'b1001000001;
  /* fppow16.vhdl:1284:24  */
  assign n4908 = x == 10'b1001000010;
  /* fppow16.vhdl:1285:24  */
  assign n4911 = x == 10'b1001000011;
  /* fppow16.vhdl:1286:24  */
  assign n4914 = x == 10'b1001000100;
  /* fppow16.vhdl:1287:24  */
  assign n4917 = x == 10'b1001000101;
  /* fppow16.vhdl:1288:24  */
  assign n4920 = x == 10'b1001000110;
  /* fppow16.vhdl:1289:24  */
  assign n4923 = x == 10'b1001000111;
  /* fppow16.vhdl:1290:24  */
  assign n4926 = x == 10'b1001001000;
  /* fppow16.vhdl:1291:24  */
  assign n4929 = x == 10'b1001001001;
  /* fppow16.vhdl:1292:24  */
  assign n4932 = x == 10'b1001001010;
  /* fppow16.vhdl:1293:24  */
  assign n4935 = x == 10'b1001001011;
  /* fppow16.vhdl:1294:24  */
  assign n4938 = x == 10'b1001001100;
  /* fppow16.vhdl:1295:24  */
  assign n4941 = x == 10'b1001001101;
  /* fppow16.vhdl:1296:24  */
  assign n4944 = x == 10'b1001001110;
  /* fppow16.vhdl:1297:24  */
  assign n4947 = x == 10'b1001001111;
  /* fppow16.vhdl:1298:24  */
  assign n4950 = x == 10'b1001010000;
  /* fppow16.vhdl:1299:24  */
  assign n4953 = x == 10'b1001010001;
  /* fppow16.vhdl:1300:24  */
  assign n4956 = x == 10'b1001010010;
  /* fppow16.vhdl:1301:24  */
  assign n4959 = x == 10'b1001010011;
  /* fppow16.vhdl:1302:24  */
  assign n4962 = x == 10'b1001010100;
  /* fppow16.vhdl:1303:24  */
  assign n4965 = x == 10'b1001010101;
  /* fppow16.vhdl:1304:24  */
  assign n4968 = x == 10'b1001010110;
  /* fppow16.vhdl:1305:24  */
  assign n4971 = x == 10'b1001010111;
  /* fppow16.vhdl:1306:24  */
  assign n4974 = x == 10'b1001011000;
  /* fppow16.vhdl:1307:24  */
  assign n4977 = x == 10'b1001011001;
  /* fppow16.vhdl:1308:24  */
  assign n4980 = x == 10'b1001011010;
  /* fppow16.vhdl:1309:24  */
  assign n4983 = x == 10'b1001011011;
  /* fppow16.vhdl:1310:24  */
  assign n4986 = x == 10'b1001011100;
  /* fppow16.vhdl:1311:24  */
  assign n4989 = x == 10'b1001011101;
  /* fppow16.vhdl:1312:24  */
  assign n4992 = x == 10'b1001011110;
  /* fppow16.vhdl:1313:24  */
  assign n4995 = x == 10'b1001011111;
  /* fppow16.vhdl:1314:24  */
  assign n4998 = x == 10'b1001100000;
  /* fppow16.vhdl:1315:24  */
  assign n5001 = x == 10'b1001100001;
  /* fppow16.vhdl:1316:24  */
  assign n5004 = x == 10'b1001100010;
  /* fppow16.vhdl:1317:24  */
  assign n5007 = x == 10'b1001100011;
  /* fppow16.vhdl:1318:24  */
  assign n5010 = x == 10'b1001100100;
  /* fppow16.vhdl:1319:24  */
  assign n5013 = x == 10'b1001100101;
  /* fppow16.vhdl:1320:24  */
  assign n5016 = x == 10'b1001100110;
  /* fppow16.vhdl:1321:24  */
  assign n5019 = x == 10'b1001100111;
  /* fppow16.vhdl:1322:24  */
  assign n5022 = x == 10'b1001101000;
  /* fppow16.vhdl:1323:24  */
  assign n5025 = x == 10'b1001101001;
  /* fppow16.vhdl:1324:24  */
  assign n5028 = x == 10'b1001101010;
  /* fppow16.vhdl:1325:24  */
  assign n5031 = x == 10'b1001101011;
  /* fppow16.vhdl:1326:24  */
  assign n5034 = x == 10'b1001101100;
  /* fppow16.vhdl:1327:24  */
  assign n5037 = x == 10'b1001101101;
  /* fppow16.vhdl:1328:24  */
  assign n5040 = x == 10'b1001101110;
  /* fppow16.vhdl:1329:24  */
  assign n5043 = x == 10'b1001101111;
  /* fppow16.vhdl:1330:24  */
  assign n5046 = x == 10'b1001110000;
  /* fppow16.vhdl:1331:24  */
  assign n5049 = x == 10'b1001110001;
  /* fppow16.vhdl:1332:24  */
  assign n5052 = x == 10'b1001110010;
  /* fppow16.vhdl:1333:24  */
  assign n5055 = x == 10'b1001110011;
  /* fppow16.vhdl:1334:24  */
  assign n5058 = x == 10'b1001110100;
  /* fppow16.vhdl:1335:24  */
  assign n5061 = x == 10'b1001110101;
  /* fppow16.vhdl:1336:24  */
  assign n5064 = x == 10'b1001110110;
  /* fppow16.vhdl:1337:24  */
  assign n5067 = x == 10'b1001110111;
  /* fppow16.vhdl:1338:24  */
  assign n5070 = x == 10'b1001111000;
  /* fppow16.vhdl:1339:24  */
  assign n5073 = x == 10'b1001111001;
  /* fppow16.vhdl:1340:24  */
  assign n5076 = x == 10'b1001111010;
  /* fppow16.vhdl:1341:24  */
  assign n5079 = x == 10'b1001111011;
  /* fppow16.vhdl:1342:24  */
  assign n5082 = x == 10'b1001111100;
  /* fppow16.vhdl:1343:24  */
  assign n5085 = x == 10'b1001111101;
  /* fppow16.vhdl:1344:24  */
  assign n5088 = x == 10'b1001111110;
  /* fppow16.vhdl:1345:24  */
  assign n5091 = x == 10'b1001111111;
  /* fppow16.vhdl:1346:24  */
  assign n5094 = x == 10'b1010000000;
  /* fppow16.vhdl:1347:24  */
  assign n5097 = x == 10'b1010000001;
  /* fppow16.vhdl:1348:24  */
  assign n5100 = x == 10'b1010000010;
  /* fppow16.vhdl:1349:24  */
  assign n5103 = x == 10'b1010000011;
  /* fppow16.vhdl:1350:24  */
  assign n5106 = x == 10'b1010000100;
  /* fppow16.vhdl:1351:24  */
  assign n5109 = x == 10'b1010000101;
  /* fppow16.vhdl:1352:24  */
  assign n5112 = x == 10'b1010000110;
  /* fppow16.vhdl:1353:24  */
  assign n5115 = x == 10'b1010000111;
  /* fppow16.vhdl:1354:24  */
  assign n5118 = x == 10'b1010001000;
  /* fppow16.vhdl:1355:24  */
  assign n5121 = x == 10'b1010001001;
  /* fppow16.vhdl:1356:24  */
  assign n5124 = x == 10'b1010001010;
  /* fppow16.vhdl:1357:24  */
  assign n5127 = x == 10'b1010001011;
  /* fppow16.vhdl:1358:24  */
  assign n5130 = x == 10'b1010001100;
  /* fppow16.vhdl:1359:24  */
  assign n5133 = x == 10'b1010001101;
  /* fppow16.vhdl:1360:24  */
  assign n5136 = x == 10'b1010001110;
  /* fppow16.vhdl:1361:24  */
  assign n5139 = x == 10'b1010001111;
  /* fppow16.vhdl:1362:24  */
  assign n5142 = x == 10'b1010010000;
  /* fppow16.vhdl:1363:24  */
  assign n5145 = x == 10'b1010010001;
  /* fppow16.vhdl:1364:24  */
  assign n5148 = x == 10'b1010010010;
  /* fppow16.vhdl:1365:24  */
  assign n5151 = x == 10'b1010010011;
  /* fppow16.vhdl:1366:24  */
  assign n5154 = x == 10'b1010010100;
  /* fppow16.vhdl:1367:24  */
  assign n5157 = x == 10'b1010010101;
  /* fppow16.vhdl:1368:24  */
  assign n5160 = x == 10'b1010010110;
  /* fppow16.vhdl:1369:24  */
  assign n5163 = x == 10'b1010010111;
  /* fppow16.vhdl:1370:24  */
  assign n5166 = x == 10'b1010011000;
  /* fppow16.vhdl:1371:24  */
  assign n5169 = x == 10'b1010011001;
  /* fppow16.vhdl:1372:24  */
  assign n5172 = x == 10'b1010011010;
  /* fppow16.vhdl:1373:24  */
  assign n5175 = x == 10'b1010011011;
  /* fppow16.vhdl:1374:24  */
  assign n5178 = x == 10'b1010011100;
  /* fppow16.vhdl:1375:24  */
  assign n5181 = x == 10'b1010011101;
  /* fppow16.vhdl:1376:24  */
  assign n5184 = x == 10'b1010011110;
  /* fppow16.vhdl:1377:24  */
  assign n5187 = x == 10'b1010011111;
  /* fppow16.vhdl:1378:24  */
  assign n5190 = x == 10'b1010100000;
  /* fppow16.vhdl:1379:24  */
  assign n5193 = x == 10'b1010100001;
  /* fppow16.vhdl:1380:24  */
  assign n5196 = x == 10'b1010100010;
  /* fppow16.vhdl:1381:24  */
  assign n5199 = x == 10'b1010100011;
  /* fppow16.vhdl:1382:24  */
  assign n5202 = x == 10'b1010100100;
  /* fppow16.vhdl:1383:24  */
  assign n5205 = x == 10'b1010100101;
  /* fppow16.vhdl:1384:24  */
  assign n5208 = x == 10'b1010100110;
  /* fppow16.vhdl:1385:24  */
  assign n5211 = x == 10'b1010100111;
  /* fppow16.vhdl:1386:24  */
  assign n5214 = x == 10'b1010101000;
  /* fppow16.vhdl:1387:24  */
  assign n5217 = x == 10'b1010101001;
  /* fppow16.vhdl:1388:24  */
  assign n5220 = x == 10'b1010101010;
  /* fppow16.vhdl:1389:24  */
  assign n5223 = x == 10'b1010101011;
  /* fppow16.vhdl:1390:24  */
  assign n5226 = x == 10'b1010101100;
  /* fppow16.vhdl:1391:24  */
  assign n5229 = x == 10'b1010101101;
  /* fppow16.vhdl:1392:24  */
  assign n5232 = x == 10'b1010101110;
  /* fppow16.vhdl:1393:24  */
  assign n5235 = x == 10'b1010101111;
  /* fppow16.vhdl:1394:24  */
  assign n5238 = x == 10'b1010110000;
  /* fppow16.vhdl:1395:24  */
  assign n5241 = x == 10'b1010110001;
  /* fppow16.vhdl:1396:24  */
  assign n5244 = x == 10'b1010110010;
  /* fppow16.vhdl:1397:24  */
  assign n5247 = x == 10'b1010110011;
  /* fppow16.vhdl:1398:24  */
  assign n5250 = x == 10'b1010110100;
  /* fppow16.vhdl:1399:24  */
  assign n5253 = x == 10'b1010110101;
  /* fppow16.vhdl:1400:24  */
  assign n5256 = x == 10'b1010110110;
  /* fppow16.vhdl:1401:24  */
  assign n5259 = x == 10'b1010110111;
  /* fppow16.vhdl:1402:24  */
  assign n5262 = x == 10'b1010111000;
  /* fppow16.vhdl:1403:24  */
  assign n5265 = x == 10'b1010111001;
  /* fppow16.vhdl:1404:24  */
  assign n5268 = x == 10'b1010111010;
  /* fppow16.vhdl:1405:24  */
  assign n5271 = x == 10'b1010111011;
  /* fppow16.vhdl:1406:24  */
  assign n5274 = x == 10'b1010111100;
  /* fppow16.vhdl:1407:24  */
  assign n5277 = x == 10'b1010111101;
  /* fppow16.vhdl:1408:24  */
  assign n5280 = x == 10'b1010111110;
  /* fppow16.vhdl:1409:24  */
  assign n5283 = x == 10'b1010111111;
  /* fppow16.vhdl:1410:24  */
  assign n5286 = x == 10'b1011000000;
  /* fppow16.vhdl:1411:24  */
  assign n5289 = x == 10'b1011000001;
  /* fppow16.vhdl:1412:24  */
  assign n5292 = x == 10'b1011000010;
  /* fppow16.vhdl:1413:24  */
  assign n5295 = x == 10'b1011000011;
  /* fppow16.vhdl:1414:24  */
  assign n5298 = x == 10'b1011000100;
  /* fppow16.vhdl:1415:24  */
  assign n5301 = x == 10'b1011000101;
  /* fppow16.vhdl:1416:24  */
  assign n5304 = x == 10'b1011000110;
  /* fppow16.vhdl:1417:24  */
  assign n5307 = x == 10'b1011000111;
  /* fppow16.vhdl:1418:24  */
  assign n5310 = x == 10'b1011001000;
  /* fppow16.vhdl:1419:24  */
  assign n5313 = x == 10'b1011001001;
  /* fppow16.vhdl:1420:24  */
  assign n5316 = x == 10'b1011001010;
  /* fppow16.vhdl:1421:24  */
  assign n5319 = x == 10'b1011001011;
  /* fppow16.vhdl:1422:24  */
  assign n5322 = x == 10'b1011001100;
  /* fppow16.vhdl:1423:24  */
  assign n5325 = x == 10'b1011001101;
  /* fppow16.vhdl:1424:24  */
  assign n5328 = x == 10'b1011001110;
  /* fppow16.vhdl:1425:24  */
  assign n5331 = x == 10'b1011001111;
  /* fppow16.vhdl:1426:24  */
  assign n5334 = x == 10'b1011010000;
  /* fppow16.vhdl:1427:24  */
  assign n5337 = x == 10'b1011010001;
  /* fppow16.vhdl:1428:24  */
  assign n5340 = x == 10'b1011010010;
  /* fppow16.vhdl:1429:24  */
  assign n5343 = x == 10'b1011010011;
  /* fppow16.vhdl:1430:24  */
  assign n5346 = x == 10'b1011010100;
  /* fppow16.vhdl:1431:24  */
  assign n5349 = x == 10'b1011010101;
  /* fppow16.vhdl:1432:24  */
  assign n5352 = x == 10'b1011010110;
  /* fppow16.vhdl:1433:24  */
  assign n5355 = x == 10'b1011010111;
  /* fppow16.vhdl:1434:24  */
  assign n5358 = x == 10'b1011011000;
  /* fppow16.vhdl:1435:24  */
  assign n5361 = x == 10'b1011011001;
  /* fppow16.vhdl:1436:24  */
  assign n5364 = x == 10'b1011011010;
  /* fppow16.vhdl:1437:24  */
  assign n5367 = x == 10'b1011011011;
  /* fppow16.vhdl:1438:24  */
  assign n5370 = x == 10'b1011011100;
  /* fppow16.vhdl:1439:24  */
  assign n5373 = x == 10'b1011011101;
  /* fppow16.vhdl:1440:24  */
  assign n5376 = x == 10'b1011011110;
  /* fppow16.vhdl:1441:24  */
  assign n5379 = x == 10'b1011011111;
  /* fppow16.vhdl:1442:24  */
  assign n5382 = x == 10'b1011100000;
  /* fppow16.vhdl:1443:24  */
  assign n5385 = x == 10'b1011100001;
  /* fppow16.vhdl:1444:24  */
  assign n5388 = x == 10'b1011100010;
  /* fppow16.vhdl:1445:24  */
  assign n5391 = x == 10'b1011100011;
  /* fppow16.vhdl:1446:24  */
  assign n5394 = x == 10'b1011100100;
  /* fppow16.vhdl:1447:24  */
  assign n5397 = x == 10'b1011100101;
  /* fppow16.vhdl:1448:24  */
  assign n5400 = x == 10'b1011100110;
  /* fppow16.vhdl:1449:24  */
  assign n5403 = x == 10'b1011100111;
  /* fppow16.vhdl:1450:24  */
  assign n5406 = x == 10'b1011101000;
  /* fppow16.vhdl:1451:24  */
  assign n5409 = x == 10'b1011101001;
  /* fppow16.vhdl:1452:24  */
  assign n5412 = x == 10'b1011101010;
  /* fppow16.vhdl:1453:24  */
  assign n5415 = x == 10'b1011101011;
  /* fppow16.vhdl:1454:24  */
  assign n5418 = x == 10'b1011101100;
  /* fppow16.vhdl:1455:24  */
  assign n5421 = x == 10'b1011101101;
  /* fppow16.vhdl:1456:24  */
  assign n5424 = x == 10'b1011101110;
  /* fppow16.vhdl:1457:24  */
  assign n5427 = x == 10'b1011101111;
  /* fppow16.vhdl:1458:24  */
  assign n5430 = x == 10'b1011110000;
  /* fppow16.vhdl:1459:24  */
  assign n5433 = x == 10'b1011110001;
  /* fppow16.vhdl:1460:24  */
  assign n5436 = x == 10'b1011110010;
  /* fppow16.vhdl:1461:24  */
  assign n5439 = x == 10'b1011110011;
  /* fppow16.vhdl:1462:24  */
  assign n5442 = x == 10'b1011110100;
  /* fppow16.vhdl:1463:24  */
  assign n5445 = x == 10'b1011110101;
  /* fppow16.vhdl:1464:24  */
  assign n5448 = x == 10'b1011110110;
  /* fppow16.vhdl:1465:24  */
  assign n5451 = x == 10'b1011110111;
  /* fppow16.vhdl:1466:24  */
  assign n5454 = x == 10'b1011111000;
  /* fppow16.vhdl:1467:24  */
  assign n5457 = x == 10'b1011111001;
  /* fppow16.vhdl:1468:24  */
  assign n5460 = x == 10'b1011111010;
  /* fppow16.vhdl:1469:24  */
  assign n5463 = x == 10'b1011111011;
  /* fppow16.vhdl:1470:24  */
  assign n5466 = x == 10'b1011111100;
  /* fppow16.vhdl:1471:24  */
  assign n5469 = x == 10'b1011111101;
  /* fppow16.vhdl:1472:24  */
  assign n5472 = x == 10'b1011111110;
  /* fppow16.vhdl:1473:24  */
  assign n5475 = x == 10'b1011111111;
  /* fppow16.vhdl:1474:24  */
  assign n5478 = x == 10'b1100000000;
  /* fppow16.vhdl:1475:24  */
  assign n5481 = x == 10'b1100000001;
  /* fppow16.vhdl:1476:24  */
  assign n5484 = x == 10'b1100000010;
  /* fppow16.vhdl:1477:24  */
  assign n5487 = x == 10'b1100000011;
  /* fppow16.vhdl:1478:24  */
  assign n5490 = x == 10'b1100000100;
  /* fppow16.vhdl:1479:24  */
  assign n5493 = x == 10'b1100000101;
  /* fppow16.vhdl:1480:24  */
  assign n5496 = x == 10'b1100000110;
  /* fppow16.vhdl:1481:24  */
  assign n5499 = x == 10'b1100000111;
  /* fppow16.vhdl:1482:24  */
  assign n5502 = x == 10'b1100001000;
  /* fppow16.vhdl:1483:24  */
  assign n5505 = x == 10'b1100001001;
  /* fppow16.vhdl:1484:24  */
  assign n5508 = x == 10'b1100001010;
  /* fppow16.vhdl:1485:24  */
  assign n5511 = x == 10'b1100001011;
  /* fppow16.vhdl:1486:24  */
  assign n5514 = x == 10'b1100001100;
  /* fppow16.vhdl:1487:24  */
  assign n5517 = x == 10'b1100001101;
  /* fppow16.vhdl:1488:24  */
  assign n5520 = x == 10'b1100001110;
  /* fppow16.vhdl:1489:24  */
  assign n5523 = x == 10'b1100001111;
  /* fppow16.vhdl:1490:24  */
  assign n5526 = x == 10'b1100010000;
  /* fppow16.vhdl:1491:24  */
  assign n5529 = x == 10'b1100010001;
  /* fppow16.vhdl:1492:24  */
  assign n5532 = x == 10'b1100010010;
  /* fppow16.vhdl:1493:24  */
  assign n5535 = x == 10'b1100010011;
  /* fppow16.vhdl:1494:24  */
  assign n5538 = x == 10'b1100010100;
  /* fppow16.vhdl:1495:24  */
  assign n5541 = x == 10'b1100010101;
  /* fppow16.vhdl:1496:24  */
  assign n5544 = x == 10'b1100010110;
  /* fppow16.vhdl:1497:24  */
  assign n5547 = x == 10'b1100010111;
  /* fppow16.vhdl:1498:24  */
  assign n5550 = x == 10'b1100011000;
  /* fppow16.vhdl:1499:24  */
  assign n5553 = x == 10'b1100011001;
  /* fppow16.vhdl:1500:24  */
  assign n5556 = x == 10'b1100011010;
  /* fppow16.vhdl:1501:24  */
  assign n5559 = x == 10'b1100011011;
  /* fppow16.vhdl:1502:24  */
  assign n5562 = x == 10'b1100011100;
  /* fppow16.vhdl:1503:24  */
  assign n5565 = x == 10'b1100011101;
  /* fppow16.vhdl:1504:24  */
  assign n5568 = x == 10'b1100011110;
  /* fppow16.vhdl:1505:24  */
  assign n5571 = x == 10'b1100011111;
  /* fppow16.vhdl:1506:24  */
  assign n5574 = x == 10'b1100100000;
  /* fppow16.vhdl:1507:24  */
  assign n5577 = x == 10'b1100100001;
  /* fppow16.vhdl:1508:24  */
  assign n5580 = x == 10'b1100100010;
  /* fppow16.vhdl:1509:24  */
  assign n5583 = x == 10'b1100100011;
  /* fppow16.vhdl:1510:24  */
  assign n5586 = x == 10'b1100100100;
  /* fppow16.vhdl:1511:24  */
  assign n5589 = x == 10'b1100100101;
  /* fppow16.vhdl:1512:24  */
  assign n5592 = x == 10'b1100100110;
  /* fppow16.vhdl:1513:24  */
  assign n5595 = x == 10'b1100100111;
  /* fppow16.vhdl:1514:24  */
  assign n5598 = x == 10'b1100101000;
  /* fppow16.vhdl:1515:24  */
  assign n5601 = x == 10'b1100101001;
  /* fppow16.vhdl:1516:24  */
  assign n5604 = x == 10'b1100101010;
  /* fppow16.vhdl:1517:24  */
  assign n5607 = x == 10'b1100101011;
  /* fppow16.vhdl:1518:24  */
  assign n5610 = x == 10'b1100101100;
  /* fppow16.vhdl:1519:24  */
  assign n5613 = x == 10'b1100101101;
  /* fppow16.vhdl:1520:24  */
  assign n5616 = x == 10'b1100101110;
  /* fppow16.vhdl:1521:24  */
  assign n5619 = x == 10'b1100101111;
  /* fppow16.vhdl:1522:24  */
  assign n5622 = x == 10'b1100110000;
  /* fppow16.vhdl:1523:24  */
  assign n5625 = x == 10'b1100110001;
  /* fppow16.vhdl:1524:24  */
  assign n5628 = x == 10'b1100110010;
  /* fppow16.vhdl:1525:24  */
  assign n5631 = x == 10'b1100110011;
  /* fppow16.vhdl:1526:24  */
  assign n5634 = x == 10'b1100110100;
  /* fppow16.vhdl:1527:24  */
  assign n5637 = x == 10'b1100110101;
  /* fppow16.vhdl:1528:24  */
  assign n5640 = x == 10'b1100110110;
  /* fppow16.vhdl:1529:24  */
  assign n5643 = x == 10'b1100110111;
  /* fppow16.vhdl:1530:24  */
  assign n5646 = x == 10'b1100111000;
  /* fppow16.vhdl:1531:24  */
  assign n5649 = x == 10'b1100111001;
  /* fppow16.vhdl:1532:24  */
  assign n5652 = x == 10'b1100111010;
  /* fppow16.vhdl:1533:24  */
  assign n5655 = x == 10'b1100111011;
  /* fppow16.vhdl:1534:24  */
  assign n5658 = x == 10'b1100111100;
  /* fppow16.vhdl:1535:24  */
  assign n5661 = x == 10'b1100111101;
  /* fppow16.vhdl:1536:24  */
  assign n5664 = x == 10'b1100111110;
  /* fppow16.vhdl:1537:24  */
  assign n5667 = x == 10'b1100111111;
  /* fppow16.vhdl:1538:24  */
  assign n5670 = x == 10'b1101000000;
  /* fppow16.vhdl:1539:24  */
  assign n5673 = x == 10'b1101000001;
  /* fppow16.vhdl:1540:24  */
  assign n5676 = x == 10'b1101000010;
  /* fppow16.vhdl:1541:24  */
  assign n5679 = x == 10'b1101000011;
  /* fppow16.vhdl:1542:24  */
  assign n5682 = x == 10'b1101000100;
  /* fppow16.vhdl:1543:24  */
  assign n5685 = x == 10'b1101000101;
  /* fppow16.vhdl:1544:24  */
  assign n5688 = x == 10'b1101000110;
  /* fppow16.vhdl:1545:24  */
  assign n5691 = x == 10'b1101000111;
  /* fppow16.vhdl:1546:24  */
  assign n5694 = x == 10'b1101001000;
  /* fppow16.vhdl:1547:24  */
  assign n5697 = x == 10'b1101001001;
  /* fppow16.vhdl:1548:24  */
  assign n5700 = x == 10'b1101001010;
  /* fppow16.vhdl:1549:24  */
  assign n5703 = x == 10'b1101001011;
  /* fppow16.vhdl:1550:24  */
  assign n5706 = x == 10'b1101001100;
  /* fppow16.vhdl:1551:24  */
  assign n5709 = x == 10'b1101001101;
  /* fppow16.vhdl:1552:24  */
  assign n5712 = x == 10'b1101001110;
  /* fppow16.vhdl:1553:24  */
  assign n5715 = x == 10'b1101001111;
  /* fppow16.vhdl:1554:24  */
  assign n5718 = x == 10'b1101010000;
  /* fppow16.vhdl:1555:24  */
  assign n5721 = x == 10'b1101010001;
  /* fppow16.vhdl:1556:24  */
  assign n5724 = x == 10'b1101010010;
  /* fppow16.vhdl:1557:24  */
  assign n5727 = x == 10'b1101010011;
  /* fppow16.vhdl:1558:24  */
  assign n5730 = x == 10'b1101010100;
  /* fppow16.vhdl:1559:24  */
  assign n5733 = x == 10'b1101010101;
  /* fppow16.vhdl:1560:24  */
  assign n5736 = x == 10'b1101010110;
  /* fppow16.vhdl:1561:24  */
  assign n5739 = x == 10'b1101010111;
  /* fppow16.vhdl:1562:24  */
  assign n5742 = x == 10'b1101011000;
  /* fppow16.vhdl:1563:24  */
  assign n5745 = x == 10'b1101011001;
  /* fppow16.vhdl:1564:24  */
  assign n5748 = x == 10'b1101011010;
  /* fppow16.vhdl:1565:24  */
  assign n5751 = x == 10'b1101011011;
  /* fppow16.vhdl:1566:24  */
  assign n5754 = x == 10'b1101011100;
  /* fppow16.vhdl:1567:24  */
  assign n5757 = x == 10'b1101011101;
  /* fppow16.vhdl:1568:24  */
  assign n5760 = x == 10'b1101011110;
  /* fppow16.vhdl:1569:24  */
  assign n5763 = x == 10'b1101011111;
  /* fppow16.vhdl:1570:24  */
  assign n5766 = x == 10'b1101100000;
  /* fppow16.vhdl:1571:24  */
  assign n5769 = x == 10'b1101100001;
  /* fppow16.vhdl:1572:24  */
  assign n5772 = x == 10'b1101100010;
  /* fppow16.vhdl:1573:24  */
  assign n5775 = x == 10'b1101100011;
  /* fppow16.vhdl:1574:24  */
  assign n5778 = x == 10'b1101100100;
  /* fppow16.vhdl:1575:24  */
  assign n5781 = x == 10'b1101100101;
  /* fppow16.vhdl:1576:24  */
  assign n5784 = x == 10'b1101100110;
  /* fppow16.vhdl:1577:24  */
  assign n5787 = x == 10'b1101100111;
  /* fppow16.vhdl:1578:24  */
  assign n5790 = x == 10'b1101101000;
  /* fppow16.vhdl:1579:24  */
  assign n5793 = x == 10'b1101101001;
  /* fppow16.vhdl:1580:24  */
  assign n5796 = x == 10'b1101101010;
  /* fppow16.vhdl:1581:24  */
  assign n5799 = x == 10'b1101101011;
  /* fppow16.vhdl:1582:24  */
  assign n5802 = x == 10'b1101101100;
  /* fppow16.vhdl:1583:24  */
  assign n5805 = x == 10'b1101101101;
  /* fppow16.vhdl:1584:24  */
  assign n5808 = x == 10'b1101101110;
  /* fppow16.vhdl:1585:24  */
  assign n5811 = x == 10'b1101101111;
  /* fppow16.vhdl:1586:24  */
  assign n5814 = x == 10'b1101110000;
  /* fppow16.vhdl:1587:24  */
  assign n5817 = x == 10'b1101110001;
  /* fppow16.vhdl:1588:24  */
  assign n5820 = x == 10'b1101110010;
  /* fppow16.vhdl:1589:24  */
  assign n5823 = x == 10'b1101110011;
  /* fppow16.vhdl:1590:24  */
  assign n5826 = x == 10'b1101110100;
  /* fppow16.vhdl:1591:24  */
  assign n5829 = x == 10'b1101110101;
  /* fppow16.vhdl:1592:24  */
  assign n5832 = x == 10'b1101110110;
  /* fppow16.vhdl:1593:24  */
  assign n5835 = x == 10'b1101110111;
  /* fppow16.vhdl:1594:24  */
  assign n5838 = x == 10'b1101111000;
  /* fppow16.vhdl:1595:24  */
  assign n5841 = x == 10'b1101111001;
  /* fppow16.vhdl:1596:24  */
  assign n5844 = x == 10'b1101111010;
  /* fppow16.vhdl:1597:24  */
  assign n5847 = x == 10'b1101111011;
  /* fppow16.vhdl:1598:24  */
  assign n5850 = x == 10'b1101111100;
  /* fppow16.vhdl:1599:24  */
  assign n5853 = x == 10'b1101111101;
  /* fppow16.vhdl:1600:24  */
  assign n5856 = x == 10'b1101111110;
  /* fppow16.vhdl:1601:24  */
  assign n5859 = x == 10'b1101111111;
  /* fppow16.vhdl:1602:24  */
  assign n5862 = x == 10'b1110000000;
  /* fppow16.vhdl:1603:24  */
  assign n5865 = x == 10'b1110000001;
  /* fppow16.vhdl:1604:24  */
  assign n5868 = x == 10'b1110000010;
  /* fppow16.vhdl:1605:24  */
  assign n5871 = x == 10'b1110000011;
  /* fppow16.vhdl:1606:24  */
  assign n5874 = x == 10'b1110000100;
  /* fppow16.vhdl:1607:24  */
  assign n5877 = x == 10'b1110000101;
  /* fppow16.vhdl:1608:24  */
  assign n5880 = x == 10'b1110000110;
  /* fppow16.vhdl:1609:24  */
  assign n5883 = x == 10'b1110000111;
  /* fppow16.vhdl:1610:24  */
  assign n5886 = x == 10'b1110001000;
  /* fppow16.vhdl:1611:24  */
  assign n5889 = x == 10'b1110001001;
  /* fppow16.vhdl:1612:24  */
  assign n5892 = x == 10'b1110001010;
  /* fppow16.vhdl:1613:24  */
  assign n5895 = x == 10'b1110001011;
  /* fppow16.vhdl:1614:24  */
  assign n5898 = x == 10'b1110001100;
  /* fppow16.vhdl:1615:24  */
  assign n5901 = x == 10'b1110001101;
  /* fppow16.vhdl:1616:24  */
  assign n5904 = x == 10'b1110001110;
  /* fppow16.vhdl:1617:24  */
  assign n5907 = x == 10'b1110001111;
  /* fppow16.vhdl:1618:24  */
  assign n5910 = x == 10'b1110010000;
  /* fppow16.vhdl:1619:24  */
  assign n5913 = x == 10'b1110010001;
  /* fppow16.vhdl:1620:24  */
  assign n5916 = x == 10'b1110010010;
  /* fppow16.vhdl:1621:24  */
  assign n5919 = x == 10'b1110010011;
  /* fppow16.vhdl:1622:24  */
  assign n5922 = x == 10'b1110010100;
  /* fppow16.vhdl:1623:24  */
  assign n5925 = x == 10'b1110010101;
  /* fppow16.vhdl:1624:24  */
  assign n5928 = x == 10'b1110010110;
  /* fppow16.vhdl:1625:24  */
  assign n5931 = x == 10'b1110010111;
  /* fppow16.vhdl:1626:24  */
  assign n5934 = x == 10'b1110011000;
  /* fppow16.vhdl:1627:24  */
  assign n5937 = x == 10'b1110011001;
  /* fppow16.vhdl:1628:24  */
  assign n5940 = x == 10'b1110011010;
  /* fppow16.vhdl:1629:24  */
  assign n5943 = x == 10'b1110011011;
  /* fppow16.vhdl:1630:24  */
  assign n5946 = x == 10'b1110011100;
  /* fppow16.vhdl:1631:24  */
  assign n5949 = x == 10'b1110011101;
  /* fppow16.vhdl:1632:24  */
  assign n5952 = x == 10'b1110011110;
  /* fppow16.vhdl:1633:24  */
  assign n5955 = x == 10'b1110011111;
  /* fppow16.vhdl:1634:24  */
  assign n5958 = x == 10'b1110100000;
  /* fppow16.vhdl:1635:24  */
  assign n5961 = x == 10'b1110100001;
  /* fppow16.vhdl:1636:24  */
  assign n5964 = x == 10'b1110100010;
  /* fppow16.vhdl:1637:24  */
  assign n5967 = x == 10'b1110100011;
  /* fppow16.vhdl:1638:24  */
  assign n5970 = x == 10'b1110100100;
  /* fppow16.vhdl:1639:24  */
  assign n5973 = x == 10'b1110100101;
  /* fppow16.vhdl:1640:24  */
  assign n5976 = x == 10'b1110100110;
  /* fppow16.vhdl:1641:24  */
  assign n5979 = x == 10'b1110100111;
  /* fppow16.vhdl:1642:24  */
  assign n5982 = x == 10'b1110101000;
  /* fppow16.vhdl:1643:24  */
  assign n5985 = x == 10'b1110101001;
  /* fppow16.vhdl:1644:24  */
  assign n5988 = x == 10'b1110101010;
  /* fppow16.vhdl:1645:24  */
  assign n5991 = x == 10'b1110101011;
  /* fppow16.vhdl:1646:24  */
  assign n5994 = x == 10'b1110101100;
  /* fppow16.vhdl:1647:24  */
  assign n5997 = x == 10'b1110101101;
  /* fppow16.vhdl:1648:24  */
  assign n6000 = x == 10'b1110101110;
  /* fppow16.vhdl:1649:24  */
  assign n6003 = x == 10'b1110101111;
  /* fppow16.vhdl:1650:24  */
  assign n6006 = x == 10'b1110110000;
  /* fppow16.vhdl:1651:24  */
  assign n6009 = x == 10'b1110110001;
  /* fppow16.vhdl:1652:24  */
  assign n6012 = x == 10'b1110110010;
  /* fppow16.vhdl:1653:24  */
  assign n6015 = x == 10'b1110110011;
  /* fppow16.vhdl:1654:24  */
  assign n6018 = x == 10'b1110110100;
  /* fppow16.vhdl:1655:24  */
  assign n6021 = x == 10'b1110110101;
  /* fppow16.vhdl:1656:24  */
  assign n6024 = x == 10'b1110110110;
  /* fppow16.vhdl:1657:24  */
  assign n6027 = x == 10'b1110110111;
  /* fppow16.vhdl:1658:24  */
  assign n6030 = x == 10'b1110111000;
  /* fppow16.vhdl:1659:24  */
  assign n6033 = x == 10'b1110111001;
  /* fppow16.vhdl:1660:24  */
  assign n6036 = x == 10'b1110111010;
  /* fppow16.vhdl:1661:24  */
  assign n6039 = x == 10'b1110111011;
  /* fppow16.vhdl:1662:24  */
  assign n6042 = x == 10'b1110111100;
  /* fppow16.vhdl:1663:24  */
  assign n6045 = x == 10'b1110111101;
  /* fppow16.vhdl:1664:24  */
  assign n6048 = x == 10'b1110111110;
  /* fppow16.vhdl:1665:24  */
  assign n6051 = x == 10'b1110111111;
  /* fppow16.vhdl:1666:24  */
  assign n6054 = x == 10'b1111000000;
  /* fppow16.vhdl:1667:24  */
  assign n6057 = x == 10'b1111000001;
  /* fppow16.vhdl:1668:24  */
  assign n6060 = x == 10'b1111000010;
  /* fppow16.vhdl:1669:24  */
  assign n6063 = x == 10'b1111000011;
  /* fppow16.vhdl:1670:24  */
  assign n6066 = x == 10'b1111000100;
  /* fppow16.vhdl:1671:24  */
  assign n6069 = x == 10'b1111000101;
  /* fppow16.vhdl:1672:24  */
  assign n6072 = x == 10'b1111000110;
  /* fppow16.vhdl:1673:24  */
  assign n6075 = x == 10'b1111000111;
  /* fppow16.vhdl:1674:24  */
  assign n6078 = x == 10'b1111001000;
  /* fppow16.vhdl:1675:24  */
  assign n6081 = x == 10'b1111001001;
  /* fppow16.vhdl:1676:24  */
  assign n6084 = x == 10'b1111001010;
  /* fppow16.vhdl:1677:24  */
  assign n6087 = x == 10'b1111001011;
  /* fppow16.vhdl:1678:24  */
  assign n6090 = x == 10'b1111001100;
  /* fppow16.vhdl:1679:24  */
  assign n6093 = x == 10'b1111001101;
  /* fppow16.vhdl:1680:24  */
  assign n6096 = x == 10'b1111001110;
  /* fppow16.vhdl:1681:24  */
  assign n6099 = x == 10'b1111001111;
  /* fppow16.vhdl:1682:24  */
  assign n6102 = x == 10'b1111010000;
  /* fppow16.vhdl:1683:24  */
  assign n6105 = x == 10'b1111010001;
  /* fppow16.vhdl:1684:24  */
  assign n6108 = x == 10'b1111010010;
  /* fppow16.vhdl:1685:24  */
  assign n6111 = x == 10'b1111010011;
  /* fppow16.vhdl:1686:24  */
  assign n6114 = x == 10'b1111010100;
  /* fppow16.vhdl:1687:24  */
  assign n6117 = x == 10'b1111010101;
  /* fppow16.vhdl:1688:24  */
  assign n6120 = x == 10'b1111010110;
  /* fppow16.vhdl:1689:24  */
  assign n6123 = x == 10'b1111010111;
  /* fppow16.vhdl:1690:24  */
  assign n6126 = x == 10'b1111011000;
  /* fppow16.vhdl:1691:24  */
  assign n6129 = x == 10'b1111011001;
  /* fppow16.vhdl:1692:24  */
  assign n6132 = x == 10'b1111011010;
  /* fppow16.vhdl:1693:24  */
  assign n6135 = x == 10'b1111011011;
  /* fppow16.vhdl:1694:24  */
  assign n6138 = x == 10'b1111011100;
  /* fppow16.vhdl:1695:24  */
  assign n6141 = x == 10'b1111011101;
  /* fppow16.vhdl:1696:24  */
  assign n6144 = x == 10'b1111011110;
  /* fppow16.vhdl:1697:24  */
  assign n6147 = x == 10'b1111011111;
  /* fppow16.vhdl:1698:24  */
  assign n6150 = x == 10'b1111100000;
  /* fppow16.vhdl:1699:24  */
  assign n6153 = x == 10'b1111100001;
  /* fppow16.vhdl:1700:24  */
  assign n6156 = x == 10'b1111100010;
  /* fppow16.vhdl:1701:24  */
  assign n6159 = x == 10'b1111100011;
  /* fppow16.vhdl:1702:24  */
  assign n6162 = x == 10'b1111100100;
  /* fppow16.vhdl:1703:24  */
  assign n6165 = x == 10'b1111100101;
  /* fppow16.vhdl:1704:24  */
  assign n6168 = x == 10'b1111100110;
  /* fppow16.vhdl:1705:24  */
  assign n6171 = x == 10'b1111100111;
  /* fppow16.vhdl:1706:24  */
  assign n6174 = x == 10'b1111101000;
  /* fppow16.vhdl:1707:24  */
  assign n6177 = x == 10'b1111101001;
  /* fppow16.vhdl:1708:24  */
  assign n6180 = x == 10'b1111101010;
  /* fppow16.vhdl:1709:24  */
  assign n6183 = x == 10'b1111101011;
  /* fppow16.vhdl:1710:24  */
  assign n6186 = x == 10'b1111101100;
  /* fppow16.vhdl:1711:24  */
  assign n6189 = x == 10'b1111101101;
  /* fppow16.vhdl:1712:24  */
  assign n6192 = x == 10'b1111101110;
  /* fppow16.vhdl:1713:24  */
  assign n6195 = x == 10'b1111101111;
  /* fppow16.vhdl:1714:24  */
  assign n6198 = x == 10'b1111110000;
  /* fppow16.vhdl:1715:24  */
  assign n6201 = x == 10'b1111110001;
  /* fppow16.vhdl:1716:24  */
  assign n6204 = x == 10'b1111110010;
  /* fppow16.vhdl:1717:24  */
  assign n6207 = x == 10'b1111110011;
  /* fppow16.vhdl:1718:24  */
  assign n6210 = x == 10'b1111110100;
  /* fppow16.vhdl:1719:24  */
  assign n6213 = x == 10'b1111110101;
  /* fppow16.vhdl:1720:24  */
  assign n6216 = x == 10'b1111110110;
  /* fppow16.vhdl:1721:24  */
  assign n6219 = x == 10'b1111110111;
  /* fppow16.vhdl:1722:24  */
  assign n6222 = x == 10'b1111111000;
  /* fppow16.vhdl:1723:24  */
  assign n6225 = x == 10'b1111111001;
  /* fppow16.vhdl:1724:24  */
  assign n6228 = x == 10'b1111111010;
  /* fppow16.vhdl:1725:24  */
  assign n6231 = x == 10'b1111111011;
  /* fppow16.vhdl:1726:24  */
  assign n6234 = x == 10'b1111111100;
  /* fppow16.vhdl:1727:24  */
  assign n6237 = x == 10'b1111111101;
  /* fppow16.vhdl:1728:24  */
  assign n6240 = x == 10'b1111111110;
  /* fppow16.vhdl:1729:24  */
  assign n6243 = x == 10'b1111111111;
  assign n6245 = {n6243, n6240, n6237, n6234, n6231, n6228, n6225, n6222, n6219, n6216, n6213, n6210, n6207, n6204, n6201, n6198, n6195, n6192, n6189, n6186, n6183, n6180, n6177, n6174, n6171, n6168, n6165, n6162, n6159, n6156, n6153, n6150, n6147, n6144, n6141, n6138, n6135, n6132, n6129, n6126, n6123, n6120, n6117, n6114, n6111, n6108, n6105, n6102, n6099, n6096, n6093, n6090, n6087, n6084, n6081, n6078, n6075, n6072, n6069, n6066, n6063, n6060, n6057, n6054, n6051, n6048, n6045, n6042, n6039, n6036, n6033, n6030, n6027, n6024, n6021, n6018, n6015, n6012, n6009, n6006, n6003, n6000, n5997, n5994, n5991, n5988, n5985, n5982, n5979, n5976, n5973, n5970, n5967, n5964, n5961, n5958, n5955, n5952, n5949, n5946, n5943, n5940, n5937, n5934, n5931, n5928, n5925, n5922, n5919, n5916, n5913, n5910, n5907, n5904, n5901, n5898, n5895, n5892, n5889, n5886, n5883, n5880, n5877, n5874, n5871, n5868, n5865, n5862, n5859, n5856, n5853, n5850, n5847, n5844, n5841, n5838, n5835, n5832, n5829, n5826, n5823, n5820, n5817, n5814, n5811, n5808, n5805, n5802, n5799, n5796, n5793, n5790, n5787, n5784, n5781, n5778, n5775, n5772, n5769, n5766, n5763, n5760, n5757, n5754, n5751, n5748, n5745, n5742, n5739, n5736, n5733, n5730, n5727, n5724, n5721, n5718, n5715, n5712, n5709, n5706, n5703, n5700, n5697, n5694, n5691, n5688, n5685, n5682, n5679, n5676, n5673, n5670, n5667, n5664, n5661, n5658, n5655, n5652, n5649, n5646, n5643, n5640, n5637, n5634, n5631, n5628, n5625, n5622, n5619, n5616, n5613, n5610, n5607, n5604, n5601, n5598, n5595, n5592, n5589, n5586, n5583, n5580, n5577, n5574, n5571, n5568, n5565, n5562, n5559, n5556, n5553, n5550, n5547, n5544, n5541, n5538, n5535, n5532, n5529, n5526, n5523, n5520, n5517, n5514, n5511, n5508, n5505, n5502, n5499, n5496, n5493, n5490, n5487, n5484, n5481, n5478, n5475, n5472, n5469, n5466, n5463, n5460, n5457, n5454, n5451, n5448, n5445, n5442, n5439, n5436, n5433, n5430, n5427, n5424, n5421, n5418, n5415, n5412, n5409, n5406, n5403, n5400, n5397, n5394, n5391, n5388, n5385, n5382, n5379, n5376, n5373, n5370, n5367, n5364, n5361, n5358, n5355, n5352, n5349, n5346, n5343, n5340, n5337, n5334, n5331, n5328, n5325, n5322, n5319, n5316, n5313, n5310, n5307, n5304, n5301, n5298, n5295, n5292, n5289, n5286, n5283, n5280, n5277, n5274, n5271, n5268, n5265, n5262, n5259, n5256, n5253, n5250, n5247, n5244, n5241, n5238, n5235, n5232, n5229, n5226, n5223, n5220, n5217, n5214, n5211, n5208, n5205, n5202, n5199, n5196, n5193, n5190, n5187, n5184, n5181, n5178, n5175, n5172, n5169, n5166, n5163, n5160, n5157, n5154, n5151, n5148, n5145, n5142, n5139, n5136, n5133, n5130, n5127, n5124, n5121, n5118, n5115, n5112, n5109, n5106, n5103, n5100, n5097, n5094, n5091, n5088, n5085, n5082, n5079, n5076, n5073, n5070, n5067, n5064, n5061, n5058, n5055, n5052, n5049, n5046, n5043, n5040, n5037, n5034, n5031, n5028, n5025, n5022, n5019, n5016, n5013, n5010, n5007, n5004, n5001, n4998, n4995, n4992, n4989, n4986, n4983, n4980, n4977, n4974, n4971, n4968, n4965, n4962, n4959, n4956, n4953, n4950, n4947, n4944, n4941, n4938, n4935, n4932, n4929, n4926, n4923, n4920, n4917, n4914, n4911, n4908, n4905, n4902, n4899, n4896, n4893, n4890, n4887, n4884, n4881, n4878, n4875, n4872, n4869, n4866, n4863, n4860, n4857, n4854, n4851, n4848, n4845, n4842, n4839, n4836, n4833, n4830, n4827, n4824, n4821, n4818, n4815, n4812, n4809, n4806, n4803, n4800, n4797, n4794, n4791, n4788, n4785, n4782, n4779, n4776, n4773, n4770, n4767, n4764, n4761, n4758, n4755, n4752, n4749, n4746, n4743, n4740, n4737, n4734, n4731, n4728, n4725, n4722, n4719, n4716, n4713, n4710, n4707, n4704, n4701, n4698, n4695, n4692, n4689, n4686, n4683, n4680, n4677, n4674, n4671, n4668, n4665, n4662, n4659, n4656, n4653, n4650, n4647, n4644, n4641, n4638, n4635, n4632, n4629, n4626, n4623, n4620, n4617, n4614, n4611, n4608, n4605, n4602, n4599, n4596, n4593, n4590, n4587, n4584, n4581, n4578, n4575, n4572, n4569, n4566, n4563, n4560, n4557, n4554, n4551, n4548, n4545, n4542, n4539, n4536, n4533, n4530, n4527, n4524, n4521, n4518, n4515, n4512, n4509, n4506, n4503, n4500, n4497, n4494, n4491, n4488, n4485, n4482, n4479, n4476, n4473, n4470, n4467, n4464, n4461, n4458, n4455, n4452, n4449, n4446, n4443, n4440, n4437, n4434, n4431, n4428, n4425, n4422, n4419, n4416, n4413, n4410, n4407, n4404, n4401, n4398, n4395, n4392, n4389, n4386, n4383, n4380, n4377, n4374, n4371, n4368, n4365, n4362, n4359, n4356, n4353, n4350, n4347, n4344, n4341, n4338, n4335, n4332, n4329, n4326, n4323, n4320, n4317, n4314, n4311, n4308, n4305, n4302, n4299, n4296, n4293, n4290, n4287, n4284, n4281, n4278, n4275, n4272, n4269, n4266, n4263, n4260, n4257, n4254, n4251, n4248, n4245, n4242, n4239, n4236, n4233, n4230, n4227, n4224, n4221, n4218, n4215, n4212, n4209, n4206, n4203, n4200, n4197, n4194, n4191, n4188, n4185, n4182, n4179, n4176, n4173, n4170, n4167, n4164, n4161, n4158, n4155, n4152, n4149, n4146, n4143, n4140, n4137, n4134, n4131, n4128, n4125, n4122, n4119, n4116, n4113, n4110, n4107, n4104, n4101, n4098, n4095, n4092, n4089, n4086, n4083, n4080, n4077, n4074, n4071, n4068, n4065, n4062, n4059, n4056, n4053, n4050, n4047, n4044, n4041, n4038, n4035, n4032, n4029, n4026, n4023, n4020, n4017, n4014, n4011, n4008, n4005, n4002, n3999, n3996, n3993, n3990, n3987, n3984, n3981, n3978, n3975, n3972, n3969, n3966, n3963, n3960, n3957, n3954, n3951, n3948, n3945, n3942, n3939, n3936, n3933, n3930, n3927, n3924, n3921, n3918, n3915, n3912, n3909, n3906, n3903, n3900, n3897, n3894, n3891, n3888, n3885, n3882, n3879, n3876, n3873, n3870, n3867, n3864, n3861, n3858, n3855, n3852, n3849, n3846, n3843, n3840, n3837, n3834, n3831, n3828, n3825, n3822, n3819, n3816, n3813, n3810, n3807, n3804, n3801, n3798, n3795, n3792, n3789, n3786, n3783, n3780, n3777, n3774, n3771, n3768, n3765, n3762, n3759, n3756, n3753, n3750, n3747, n3744, n3741, n3738, n3735, n3732, n3729, n3726, n3723, n3720, n3717, n3714, n3711, n3708, n3705, n3702, n3699, n3696, n3693, n3690, n3687, n3684, n3681, n3678, n3675, n3672, n3669, n3666, n3663, n3660, n3657, n3654, n3651, n3648, n3645, n3642, n3639, n3636, n3633, n3630, n3627, n3624, n3621, n3618, n3615, n3612, n3609, n3606, n3603, n3600, n3597, n3594, n3591, n3588, n3585, n3582, n3579, n3576, n3573, n3570, n3567, n3564, n3561, n3558, n3555, n3552, n3549, n3546, n3543, n3540, n3537, n3534, n3531, n3528, n3525, n3522, n3519, n3516, n3513, n3510, n3507, n3504, n3501, n3498, n3495, n3492, n3489, n3486, n3483, n3480, n3477, n3474, n3471, n3468, n3465, n3462, n3459, n3456, n3453, n3450, n3447, n3444, n3441, n3438, n3435, n3432, n3429, n3426, n3423, n3420, n3417, n3414, n3411, n3408, n3405, n3402, n3399, n3396, n3393, n3390, n3387, n3384, n3381, n3378, n3375, n3372, n3369, n3366, n3363, n3360, n3357, n3354, n3351, n3348, n3345, n3342, n3339, n3336, n3333, n3330, n3327, n3324, n3321, n3318, n3315, n3312, n3309, n3306, n3303, n3300, n3297, n3294, n3291, n3288, n3285, n3282, n3279, n3276, n3273, n3270, n3267, n3264, n3261, n3258, n3255, n3252, n3249, n3246, n3243, n3240, n3237, n3234, n3231, n3228, n3225, n3222, n3219, n3216, n3213, n3210, n3207, n3204, n3201, n3198, n3195, n3192, n3189, n3186, n3183, n3180, n3177, n3174};
  /* fppow16.vhdl:705:4  */
  always @*
    case (n6245)
      1024'b1000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01111111111000;
      1024'b0100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01111111110000;
      1024'b0010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01111111101000;
      1024'b0001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01111111100000;
      1024'b0000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01111111011000;
      1024'b0000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01111111010000;
      1024'b0000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01111111001000;
      1024'b0000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01111111000000;
      1024'b0000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01111110111000;
      1024'b0000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01111110110000;
      1024'b0000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01111110101000;
      1024'b0000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01111110100001;
      1024'b0000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01111110011001;
      1024'b0000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01111110010001;
      1024'b0000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01111110001001;
      1024'b0000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01111110000001;
      1024'b0000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01111101111001;
      1024'b0000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01111101110001;
      1024'b0000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01111101101001;
      1024'b0000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01111101100010;
      1024'b0000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01111101011010;
      1024'b0000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01111101010010;
      1024'b0000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01111101001010;
      1024'b0000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01111101000010;
      1024'b0000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01111100111010;
      1024'b0000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01111100110011;
      1024'b0000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01111100101011;
      1024'b0000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01111100100011;
      1024'b0000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01111100011011;
      1024'b0000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01111100010011;
      1024'b0000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01111100001100;
      1024'b0000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01111100000100;
      1024'b0000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01111011111100;
      1024'b0000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01111011110100;
      1024'b0000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01111011101101;
      1024'b0000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01111011100101;
      1024'b0000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01111011011101;
      1024'b0000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01111011010110;
      1024'b0000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01111011001110;
      1024'b0000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01111011000110;
      1024'b0000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01111010111110;
      1024'b0000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01111010110111;
      1024'b0000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01111010101111;
      1024'b0000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01111010100111;
      1024'b0000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01111010100000;
      1024'b0000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01111010011000;
      1024'b0000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01111010010000;
      1024'b0000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01111010001001;
      1024'b0000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01111010000001;
      1024'b0000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01111001111010;
      1024'b0000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01111001110010;
      1024'b0000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01111001101010;
      1024'b0000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01111001100011;
      1024'b0000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01111001011011;
      1024'b0000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01111001010100;
      1024'b0000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01111001001100;
      1024'b0000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01111001000100;
      1024'b0000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01111000111101;
      1024'b0000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01111000110101;
      1024'b0000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01111000101110;
      1024'b0000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01111000100110;
      1024'b0000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01111000011111;
      1024'b0000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01111000010111;
      1024'b0000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01111000010000;
      1024'b0000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01111000001000;
      1024'b0000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01111000000001;
      1024'b0000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01110111111001;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01110111110010;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01110111101010;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01110111100011;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01110111011011;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01110111010100;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01110111001100;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01110111000101;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01110110111101;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01110110110110;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01110110101111;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01110110100111;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01110110100000;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01110110011000;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01110110010001;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01110110001010;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01110110000010;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01110101111011;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01110101110011;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01110101101100;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01110101100101;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01110101011101;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01110101010110;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01110101001111;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01110101000111;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01110101000000;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01110100111001;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01110100110001;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01110100101010;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01110100100011;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01110100011100;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01110100010100;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01110100001101;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01110100000110;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01110011111111;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01110011110111;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01110011110000;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01110011101001;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01110011100010;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01110011011010;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01110011010011;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01110011001100;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01110011000101;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01110010111110;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01110010110110;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01110010101111;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01110010101000;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01110010100001;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01110010011010;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01110010010011;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01110010001011;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01110010000100;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01110001111101;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01110001110110;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01110001101111;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01110001101000;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01110001100001;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01110001011010;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01110001010011;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01110001001100;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01110001000100;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01110000111101;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01110000110110;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01110000101111;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01110000101000;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01110000100001;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01110000011010;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01110000010011;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01110000001100;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01110000000101;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01101111111110;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01101111110111;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01101111110000;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01101111101001;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01101111100010;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01101111011011;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01101111010100;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01101111001101;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01101111000110;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01101110111111;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01101110111001;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01101110110010;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01101110101011;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01101110100100;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01101110011101;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01101110010110;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01101110001111;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01101110001000;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01101110000001;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01101101111010;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01101101110100;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01101101101101;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01101101100110;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01101101011111;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01101101011000;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01101101010001;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01101101001010;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01101101000100;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01101100111101;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01101100110110;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01101100101111;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01101100101000;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01101100100010;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01101100011011;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01101100010100;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01101100001101;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01101100000111;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01101100000000;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01101011111001;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01101011110010;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01101011101100;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01101011100101;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01101011011110;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01101011010111;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01101011010001;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01101011001010;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01101011000011;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01101010111101;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01101010110110;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01101010101111;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01101010101001;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01101010100010;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01101010011011;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01101010010101;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01101010001110;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01101010000111;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01101010000001;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01101001111010;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01101001110100;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01101001101101;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01101001100110;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01101001100000;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01101001011001;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01101001010011;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01101001001100;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01101001000101;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01101000111111;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01101000111000;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01101000110010;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01101000101011;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01101000100101;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01101000011110;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01101000011000;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01101000010001;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01101000001011;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01101000000100;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01100111111110;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01100111110111;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01100111110001;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01100111101010;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01100111100100;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01100111011101;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01100111010111;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01100111010000;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01100111001010;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01100111000011;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01100110111101;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01100110110110;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01100110110000;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01100110101010;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01100110100011;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01100110011101;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01100110010110;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01100110010000;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01100110001010;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01100110000011;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01100101111101;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01100101110110;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01100101110000;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01100101101010;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01100101100011;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01100101011101;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01100101010111;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01100101010000;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01100101001010;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01100101000100;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01100100111101;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01100100110111;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01100100110001;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01100100101011;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01100100100100;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01100100011110;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01100100011000;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01100100010001;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01100100001011;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01100100000101;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01100011111111;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01100011111000;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01100011110010;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01100011101100;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01100011100110;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01100011011111;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01100011011001;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01100011010011;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01100011001101;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01100011000111;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01100011000000;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01100010111010;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01100010110100;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01100010101110;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01100010101000;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01100010100010;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01100010011011;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01100010010101;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01100010001111;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01100010001001;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01100010000011;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01100001111101;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01100001110111;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01100001110001;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01100001101010;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01100001100100;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01100001011110;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01100001011000;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01100001010010;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01100001001100;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01100001000110;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01100001000000;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01100000111010;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01100000110100;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01100000101110;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01100000101000;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01100000100010;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01100000011100;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01100000010110;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01100000010000;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01100000001010;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01100000000100;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01011111111110;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01011111111000;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01011111110010;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01011111101100;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01011111100110;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01011111100000;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01011111011010;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01011111010100;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01011111001110;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01011111001000;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01011111000010;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01011110111100;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01011110110110;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01011110110000;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01011110101010;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01011110100100;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01011110011110;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01011110011000;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01011110010011;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01011110001101;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01011110000111;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01011110000001;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01011101111011;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01011101110101;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01011101101111;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01011101101001;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01011101100100;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01011101011110;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01011101011000;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01011101010010;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01011101001100;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01011101000110;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01011101000001;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01011100111011;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01011100110101;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01011100101111;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01011100101001;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01011100100100;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01011100011110;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01011100011000;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01011100010010;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01011100001100;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01011100000111;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01011100000001;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01011011111011;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01011011110101;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01011011110000;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01011011101010;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01011011100100;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01011011011111;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01011011011001;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01011011010011;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01011011001101;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01011011001000;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01011011000010;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01011010111100;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01011010110111;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01011010110001;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01011010101011;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01011010100110;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01011010100000;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01011010011010;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01011010010101;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01011010001111;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01011010001001;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01011010000100;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01011001111110;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01011001111001;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01011001110011;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01011001101101;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01011001101000;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01011001100010;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01011001011101;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01011001010111;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01011001010001;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01011001001100;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01011001000110;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01011001000001;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01011000111011;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01011000110110;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01011000110000;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01011000101010;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01011000100101;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01011000011111;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01011000011010;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01011000010100;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01011000001111;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01011000001001;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01011000000100;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01010111111110;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01010111111001;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01010111110011;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01010111101110;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01010111101000;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01010111100011;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01010111011101;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01010111011000;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01010111010010;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01010111001101;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01010111001000;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01010111000010;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01010110111101;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01010110110111;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01010110110010;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01010110101100;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01010110100111;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01010110100010;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01010110011100;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01010110010111;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01010110010001;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01010110001100;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01010110000111;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01010110000001;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01010101111100;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01010101110110;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01010101110001;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01010101101100;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01010101100110;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01010101100001;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01010101011100;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01010101010110;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01010101010001;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01010101001100;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01010101000110;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01010101000001;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01010100111100;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01010100110110;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01010100110001;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01010100101100;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01010100100111;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01010100100001;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01010100011100;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01010100010111;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01010100010001;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01010100001100;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01010100000111;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01010100000010;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01010011111100;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01010011110111;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01010011110010;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01010011101101;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01010011100111;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01010011100010;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01010011011101;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01010011011000;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01010011010011;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01010011001101;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01010011001000;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01010011000011;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01010010111110;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01010010111001;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01010010110011;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01010010101110;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01010010101001;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01010010100100;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01010010011111;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01010010011010;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01010010010101;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01010010001111;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01010010001010;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01010010000101;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01010010000000;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01010001111011;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01010001110110;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01010001110001;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01010001101100;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01010001100110;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01010001100001;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01010001011100;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01010001010111;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01010001010010;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01010001001101;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01010001001000;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01010001000011;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01010000111110;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01010000111001;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01010000110100;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01010000101111;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01010000101010;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01010000100101;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01010000100000;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01010000011010;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01010000010101;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01010000010000;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01010000001011;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01010000000110;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01010000000001;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01001111111100;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01001111110111;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01001111110010;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01001111101101;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01001111101000;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01001111100011;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01001111011111;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01001111011010;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01001111010101;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01001111010000;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01001111001011;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01001111000110;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01001111000001;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01001110111100;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01001110110111;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01001110110010;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01001110101101;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01001110101000;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01001110100011;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01001110011110;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01001110011001;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01001110010101;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01001110010000;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01001110001011;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01001110000110;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01001110000001;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01001101111100;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01001101110111;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01001101110010;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01001101101110;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b01001101101001;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b11010010110101;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b11010010101000;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b11010010011011;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b11010010001110;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b11010010000001;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b11010001110011;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b11010001100110;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b11010001011001;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b11010001001100;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b11010000111111;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b11010000110010;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b11010000100101;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b11010000011000;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b11010000001011;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b11001111111110;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b11001111110001;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b11001111100100;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b11001111010111;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b11001111001010;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b11001110111101;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b11001110110000;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b11001110100011;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b11001110010110;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b11001110001001;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b11001101111101;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b11001101110000;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b11001101100011;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b11001101010110;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b11001101001001;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b11001100111100;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b11001100110000;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b11001100100011;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b11001100010110;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b11001100001001;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b11001011111100;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b11001011110000;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b11001011100011;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b11001011010110;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b11001011001010;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b11001010111101;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b11001010110000;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b11001010100100;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b11001010010111;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b11001010001010;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b11001001111110;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b11001001110001;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b11001001100100;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b11001001011000;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b11001001001011;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b11001000111111;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b11001000110010;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b11001000100110;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b11001000011001;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b11001000001101;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b11001000000000;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b11000111110100;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b11000111100111;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b11000111011011;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b11000111001110;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b11000111000010;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b11000110110101;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b11000110101001;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b11000110011100;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b11000110010000;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b11000110000100;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b11000101110111;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b11000101101011;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b11000101011111;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b11000101010010;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b11000101000110;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b11000100111010;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b11000100101101;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b11000100100001;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b11000100010101;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b11000100001000;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b11000011111100;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b11000011110000;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b11000011100100;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b11000011011000;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b11000011001011;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b11000010111111;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b11000010110011;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b11000010100111;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b11000010011011;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b11000010001110;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b11000010000010;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b11000001110110;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b11000001101010;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b11000001011110;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b11000001010010;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b11000001000110;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b11000000111010;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b11000000101110;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b11000000100010;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b11000000010110;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b11000000001010;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b10111111111110;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b10111111110010;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b10111111100110;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b10111111011010;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b10111111001110;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b10111111000010;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b10111110110110;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b10111110101010;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b10111110011110;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b10111110010010;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b10111110000110;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b10111101111010;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b10111101101111;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b10111101100011;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b10111101010111;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b10111101001011;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b10111100111111;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b10111100110011;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b10111100101000;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b10111100011100;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b10111100010000;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b10111100000100;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b10111011111001;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b10111011101101;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b10111011100001;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b10111011010101;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b10111011001010;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b10111010111110;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b10111010110010;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b10111010100111;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b10111010011011;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b10111010001111;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b10111010000100;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b10111001111000;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b10111001101100;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b10111001100001;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b10111001010101;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b10111001001010;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b10111000111110;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b10111000110011;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b10111000100111;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b10111000011011;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b10111000010000;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b10111000000100;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b10110111111001;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b10110111101101;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b10110111100010;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b10110111010110;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b10110111001011;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b10110111000000;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b10110110110100;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b10110110101001;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b10110110011101;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b10110110010010;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b10110110000111;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b10110101111011;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b10110101110000;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b10110101100100;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b10110101011001;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b10110101001110;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b10110101000010;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b10110100110111;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b10110100101100;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b10110100100001;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b10110100010101;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b10110100001010;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b10110011111111;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b10110011110100;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b10110011101000;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b10110011011101;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b10110011010010;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b10110011000111;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b10110010111011;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b10110010110000;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b10110010100101;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b10110010011010;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b10110010001111;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b10110010000100;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b10110001111001;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b10110001101101;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b10110001100010;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b10110001010111;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b10110001001100;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b10110001000001;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b10110000110110;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b10110000101011;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b10110000100000;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b10110000010101;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b10110000001010;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b10101111111111;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b10101111110100;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b10101111101001;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b10101111011110;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b10101111010011;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b10101111001000;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b10101110111101;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b10101110110010;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b10101110100111;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b10101110011100;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b10101110010001;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b10101110000111;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b10101101111100;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b10101101110001;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b10101101100110;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b10101101011011;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b10101101010000;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b10101101000101;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b10101100111011;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b10101100110000;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b10101100100101;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b10101100011010;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b10101100010000;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b10101100000101;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b10101011111010;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b10101011101111;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b10101011100101;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b10101011011010;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b10101011001111;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b10101011000100;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b10101010111010;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b10101010101111;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b10101010100100;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b10101010011010;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b10101010001111;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b10101010000100;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b10101001111010;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b10101001101111;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b10101001100101;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b10101001011010;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b10101001001111;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b10101001000101;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b10101000111010;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b10101000110000;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b10101000100101;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b10101000011011;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b10101000010000;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b10101000000110;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b10100111111011;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b10100111110001;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b10100111100110;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b10100111011100;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b10100111010001;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b10100111000111;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b10100110111100;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b10100110110010;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b10100110101000;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b10100110011101;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b10100110010011;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b10100110001000;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b10100101111110;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b10100101110100;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b10100101101001;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b10100101011111;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b10100101010101;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b10100101001010;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b10100101000000;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b10100100110110;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b10100100101011;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b10100100100001;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b10100100010111;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b10100100001100;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b10100100000010;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b10100011111000;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b10100011101110;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b10100011100100;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b10100011011001;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b10100011001111;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b10100011000101;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b10100010111011;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b10100010110001;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b10100010100110;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b10100010011100;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b10100010010010;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b10100010001000;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b10100001111110;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b10100001110100;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b10100001101010;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b10100001011111;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b10100001010101;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b10100001001011;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b10100001000001;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b10100000110111;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b10100000101101;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b10100000100011;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b10100000011001;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b10100000001111;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b10100000000101;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b10011111111011;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b10011111110001;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b10011111100111;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b10011111011101;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b10011111010011;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b10011111001001;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b10011110111111;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b10011110110101;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b10011110101011;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b10011110100001;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b10011110011000;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b10011110001110;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b10011110000100;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b10011101111010;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b10011101110000;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b10011101100110;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b10011101011100;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b10011101010010;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b10011101001001;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b10011100111111;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b10011100110101;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b10011100101011;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b10011100100001;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b10011100011000;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b10011100001110;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b10011100000100;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b10011011111010;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b10011011110001;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b10011011100111;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b10011011011101;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b10011011010100;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b10011011001010;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b10011011000000;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b10011010110110;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b10011010101101;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b10011010100011;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b10011010011001;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b10011010010000;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b10011010000110;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b10011001111101;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b10011001110011;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b10011001101001;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b10011001100000;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b10011001010110;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b10011001001101;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b10011001000011;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b10011000111001;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b10011000110000;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b10011000100110;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b10011000011101;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b10011000010011;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b10011000001010;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b10011000000000;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b10010111110111;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b10010111101101;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b10010111100100;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b10010111011010;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b10010111010001;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b10010111000111;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b10010110111110;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b10010110110101;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b10010110101011;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b10010110100010;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b10010110011000;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b10010110001111;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b10010110000110;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b10010101111100;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b10010101110011;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b10010101101001;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b10010101100000;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b10010101010111;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b10010101001101;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b10010101000100;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b10010100111011;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b10010100110001;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b10010100101000;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b10010100011111;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b10010100010110;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b10010100001100;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b10010100000011;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b10010011111010;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b10010011110001;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b10010011100111;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b10010011011110;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b10010011010101;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b10010011001100;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b10010011000011;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b10010010111001;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b10010010110000;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b10010010100111;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b10010010011110;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b10010010010101;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b10010010001100;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b10010010000010;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b10010001111001;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b10010001110000;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b10010001100111;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b10010001011110;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b10010001010101;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b10010001001100;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b10010001000011;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b10010000111010;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b10010000110001;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b10010000101000;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b10010000011111;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b10010000010110;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b10010000001101;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b10010000000100;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b10001111111011;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b10001111110010;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b10001111101001;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b10001111100000;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b10001111010111;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b10001111001110;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b10001111000101;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b10001110111100;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b10001110110011;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b10001110101010;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b10001110100001;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b10001110011000;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b10001110001111;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b10001110000110;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b10001101111101;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b10001101110101;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b10001101101100;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b10001101100011;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b10001101011010;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b10001101010001;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b10001101001000;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b10001101000000;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b10001100110111;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b10001100101110;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b10001100100101;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b10001100011100;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b10001100010100;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b10001100001011;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b10001100000010;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b10001011111001;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b10001011110001;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b10001011101000;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b10001011011111;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b10001011010110;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b10001011001110;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b10001011000101;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b10001010111100;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b10001010110100;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b10001010101011;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b10001010100010;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b10001010011010;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b10001010010001;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b10001010001000;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b10001010000000;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b10001001110111;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b10001001101111;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b10001001100110;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b10001001011101;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b10001001010101;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b10001001001100;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b10001001000100;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b10001000111011;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b10001000110010;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b10001000101010;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b10001000100001;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b10001000011001;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b10001000010000;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b10001000001000;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b10000111111111;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b10000111110111;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000: n6246 = 14'b10000111101110;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000: n6246 = 14'b10000111100110;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000: n6246 = 14'b10000111011101;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000: n6246 = 14'b10000111010101;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000: n6246 = 14'b10000111001100;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000: n6246 = 14'b10000111000100;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000: n6246 = 14'b10000110111100;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000: n6246 = 14'b10000110110011;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000: n6246 = 14'b10000110101011;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000: n6246 = 14'b10000110100010;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000: n6246 = 14'b10000110011010;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000: n6246 = 14'b10000110010010;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000: n6246 = 14'b10000110001001;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000: n6246 = 14'b10000110000001;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000: n6246 = 14'b10000101111000;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000: n6246 = 14'b10000101110000;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000: n6246 = 14'b10000101101000;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000: n6246 = 14'b10000101011111;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000: n6246 = 14'b10000101010111;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000: n6246 = 14'b10000101001111;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000: n6246 = 14'b10000101000110;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000: n6246 = 14'b10000100111110;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000: n6246 = 14'b10000100110110;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000: n6246 = 14'b10000100101101;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000: n6246 = 14'b10000100100101;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000: n6246 = 14'b10000100011101;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000: n6246 = 14'b10000100010101;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000: n6246 = 14'b10000100001100;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000: n6246 = 14'b10000100000100;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000: n6246 = 14'b10000011111100;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000: n6246 = 14'b10000011110100;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000: n6246 = 14'b10000011101011;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000: n6246 = 14'b10000011100011;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000: n6246 = 14'b10000011011011;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000: n6246 = 14'b10000011010011;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000: n6246 = 14'b10000011001010;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000: n6246 = 14'b10000011000010;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000: n6246 = 14'b10000010111010;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000: n6246 = 14'b10000010110010;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000: n6246 = 14'b10000010101010;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000: n6246 = 14'b10000010100010;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000: n6246 = 14'b10000010011001;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000: n6246 = 14'b10000010010001;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000: n6246 = 14'b10000010001001;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000: n6246 = 14'b10000010000001;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000: n6246 = 14'b10000001111001;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000: n6246 = 14'b10000001110001;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000: n6246 = 14'b10000001101001;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000: n6246 = 14'b10000001100001;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000: n6246 = 14'b10000001011000;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000: n6246 = 14'b10000001010000;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000: n6246 = 14'b10000001001000;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000: n6246 = 14'b10000001000000;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000: n6246 = 14'b10000000111000;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000: n6246 = 14'b10000000110000;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000: n6246 = 14'b10000000101000;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000: n6246 = 14'b10000000100000;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000: n6246 = 14'b10000000011000;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100: n6246 = 14'b10000000010000;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010: n6246 = 14'b10000000001000;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001: n6246 = 14'b10000000000000;
      default: n6246 = 14'bX;
    endcase
endmodule

module intadder_13_freq500_uid92
  (input  clk,
   input  [12:0] x,
   input  [12:0] y,
   input  cin,
   output [12:0] r);
  wire [12:0] rtmp;
  wire [12:0] x_d1;
  wire [12:0] x_d2;
  wire [12:0] y_d1;
  wire cin_d1;
  wire cin_d2;
  wire cin_d3;
  wire cin_d4;
  wire cin_d5;
  wire cin_d6;
  wire cin_d7;
  wire cin_d8;
  wire cin_d9;
  wire cin_d10;
  wire cin_d11;
  wire cin_d12;
  wire cin_d13;
  wire cin_d14;
  wire cin_d15;
  wire cin_d16;
  wire [12:0] n3149;
  wire [12:0] n3150;
  wire [12:0] n3151;
  reg [12:0] n3152;
  reg [12:0] n3153;
  reg [12:0] n3154;
  reg n3155;
  reg n3156;
  reg n3157;
  reg n3158;
  reg n3159;
  reg n3160;
  reg n3161;
  reg n3162;
  reg n3163;
  reg n3164;
  reg n3165;
  reg n3166;
  reg n3167;
  reg n3168;
  reg n3169;
  reg n3170;
  assign r = rtmp; //(module output)
  /* fppow16.vhdl:4112:8  */
  assign rtmp = n3151; // (signal)
  /* fppow16.vhdl:4114:8  */
  assign x_d1 = n3152; // (signal)
  /* fppow16.vhdl:4114:14  */
  assign x_d2 = n3153; // (signal)
  /* fppow16.vhdl:4116:8  */
  assign y_d1 = n3154; // (signal)
  /* fppow16.vhdl:4118:8  */
  assign cin_d1 = n3155; // (signal)
  /* fppow16.vhdl:4118:16  */
  assign cin_d2 = n3156; // (signal)
  /* fppow16.vhdl:4118:24  */
  assign cin_d3 = n3157; // (signal)
  /* fppow16.vhdl:4118:32  */
  assign cin_d4 = n3158; // (signal)
  /* fppow16.vhdl:4118:40  */
  assign cin_d5 = n3159; // (signal)
  /* fppow16.vhdl:4118:48  */
  assign cin_d6 = n3160; // (signal)
  /* fppow16.vhdl:4118:56  */
  assign cin_d7 = n3161; // (signal)
  /* fppow16.vhdl:4118:64  */
  assign cin_d8 = n3162; // (signal)
  /* fppow16.vhdl:4118:72  */
  assign cin_d9 = n3163; // (signal)
  /* fppow16.vhdl:4118:80  */
  assign cin_d10 = n3164; // (signal)
  /* fppow16.vhdl:4118:89  */
  assign cin_d11 = n3165; // (signal)
  /* fppow16.vhdl:4118:98  */
  assign cin_d12 = n3166; // (signal)
  /* fppow16.vhdl:4118:107  */
  assign cin_d13 = n3167; // (signal)
  /* fppow16.vhdl:4118:116  */
  assign cin_d14 = n3168; // (signal)
  /* fppow16.vhdl:4118:125  */
  assign cin_d15 = n3169; // (signal)
  /* fppow16.vhdl:4118:134  */
  assign cin_d16 = n3170; // (signal)
  /* fppow16.vhdl:4145:17  */
  assign n3149 = x_d2 + y_d1;
  /* fppow16.vhdl:4145:24  */
  assign n3150 = {12'b0, cin_d16};  //  uext
  /* fppow16.vhdl:4145:24  */
  assign n3151 = n3149 + n3150;
  /* fppow16.vhdl:4123:10  */
  always @(posedge clk)
    n3152 <= x;
  /* fppow16.vhdl:4123:10  */
  always @(posedge clk)
    n3153 <= x_d1;
  /* fppow16.vhdl:4123:10  */
  always @(posedge clk)
    n3154 <= y;
  /* fppow16.vhdl:4123:10  */
  always @(posedge clk)
    n3155 <= cin;
  /* fppow16.vhdl:4123:10  */
  always @(posedge clk)
    n3156 <= cin_d1;
  /* fppow16.vhdl:4123:10  */
  always @(posedge clk)
    n3157 <= cin_d2;
  /* fppow16.vhdl:4123:10  */
  always @(posedge clk)
    n3158 <= cin_d3;
  /* fppow16.vhdl:4123:10  */
  always @(posedge clk)
    n3159 <= cin_d4;
  /* fppow16.vhdl:4123:10  */
  always @(posedge clk)
    n3160 <= cin_d5;
  /* fppow16.vhdl:4123:10  */
  always @(posedge clk)
    n3161 <= cin_d6;
  /* fppow16.vhdl:4123:10  */
  always @(posedge clk)
    n3162 <= cin_d7;
  /* fppow16.vhdl:4123:10  */
  always @(posedge clk)
    n3163 <= cin_d8;
  /* fppow16.vhdl:4123:10  */
  always @(posedge clk)
    n3164 <= cin_d9;
  /* fppow16.vhdl:4123:10  */
  always @(posedge clk)
    n3165 <= cin_d10;
  /* fppow16.vhdl:4123:10  */
  always @(posedge clk)
    n3166 <= cin_d11;
  /* fppow16.vhdl:4123:10  */
  always @(posedge clk)
    n3167 <= cin_d12;
  /* fppow16.vhdl:4123:10  */
  always @(posedge clk)
    n3168 <= cin_d13;
  /* fppow16.vhdl:4123:10  */
  always @(posedge clk)
    n3169 <= cin_d14;
  /* fppow16.vhdl:4123:10  */
  always @(posedge clk)
    n3170 <= cin_d15;
endmodule

module fixrealkcm_freq500_uid84
  (input  clk,
   input  [4:0] x,
   output [17:0] r);
  wire [4:0] fixrealkcm_freq500_uid84_a0;
  wire [17:0] fixrealkcm_freq500_uid84_t0;
  wire [17:0] fixrealkcm_freq500_uid84_t0_copy88;
  wire bh85_w0_0;
  wire bh85_w1_0;
  wire bh85_w2_0;
  wire bh85_w3_0;
  wire bh85_w4_0;
  wire bh85_w5_0;
  wire bh85_w6_0;
  wire bh85_w7_0;
  wire bh85_w8_0;
  wire bh85_w9_0;
  wire bh85_w10_0;
  wire bh85_w11_0;
  wire bh85_w12_0;
  wire bh85_w13_0;
  wire bh85_w14_0;
  wire bh85_w15_0;
  wire bh85_w16_0;
  wire bh85_w17_0;
  wire [17:0] tmp_bitheapresult_bh85_17;
  wire [17:0] bitheapresult_bh85;
  wire [17:0] outres;
  wire [17:0] fixrealkcm_freq500_uid84_table0_n3087;
  wire n3090;
  wire n3091;
  wire n3092;
  wire n3093;
  wire n3094;
  wire n3095;
  wire n3096;
  wire n3097;
  wire n3098;
  wire n3099;
  wire n3100;
  wire n3101;
  wire n3102;
  wire n3103;
  wire n3104;
  wire n3105;
  wire n3106;
  wire n3107;
  wire [1:0] n3108;
  wire [2:0] n3109;
  wire [3:0] n3110;
  wire [4:0] n3111;
  wire [5:0] n3112;
  wire [6:0] n3113;
  wire [7:0] n3114;
  wire [8:0] n3115;
  wire [9:0] n3116;
  wire [10:0] n3117;
  wire [11:0] n3118;
  wire [12:0] n3119;
  wire [13:0] n3120;
  wire [14:0] n3121;
  wire [15:0] n3122;
  wire [16:0] n3123;
  wire [17:0] n3124;
  assign r = outres; //(module output)
  /* fppow16.vhdl:3999:8  */
  assign fixrealkcm_freq500_uid84_t0 = fixrealkcm_freq500_uid84_t0_copy88; // (signal)
  /* fppow16.vhdl:4001:8  */
  assign fixrealkcm_freq500_uid84_t0_copy88 = fixrealkcm_freq500_uid84_table0_n3087; // (signal)
  /* fppow16.vhdl:4003:8  */
  assign bh85_w0_0 = n3090; // (signal)
  /* fppow16.vhdl:4005:8  */
  assign bh85_w1_0 = n3091; // (signal)
  /* fppow16.vhdl:4007:8  */
  assign bh85_w2_0 = n3092; // (signal)
  /* fppow16.vhdl:4009:8  */
  assign bh85_w3_0 = n3093; // (signal)
  /* fppow16.vhdl:4011:8  */
  assign bh85_w4_0 = n3094; // (signal)
  /* fppow16.vhdl:4013:8  */
  assign bh85_w5_0 = n3095; // (signal)
  /* fppow16.vhdl:4015:8  */
  assign bh85_w6_0 = n3096; // (signal)
  /* fppow16.vhdl:4017:8  */
  assign bh85_w7_0 = n3097; // (signal)
  /* fppow16.vhdl:4019:8  */
  assign bh85_w8_0 = n3098; // (signal)
  /* fppow16.vhdl:4021:8  */
  assign bh85_w9_0 = n3099; // (signal)
  /* fppow16.vhdl:4023:8  */
  assign bh85_w10_0 = n3100; // (signal)
  /* fppow16.vhdl:4025:8  */
  assign bh85_w11_0 = n3101; // (signal)
  /* fppow16.vhdl:4027:8  */
  assign bh85_w12_0 = n3102; // (signal)
  /* fppow16.vhdl:4029:8  */
  assign bh85_w13_0 = n3103; // (signal)
  /* fppow16.vhdl:4031:8  */
  assign bh85_w14_0 = n3104; // (signal)
  /* fppow16.vhdl:4033:8  */
  assign bh85_w15_0 = n3105; // (signal)
  /* fppow16.vhdl:4035:8  */
  assign bh85_w16_0 = n3106; // (signal)
  /* fppow16.vhdl:4037:8  */
  assign bh85_w17_0 = n3107; // (signal)
  /* fppow16.vhdl:4039:8  */
  assign tmp_bitheapresult_bh85_17 = n3124; // (signal)
  /* fppow16.vhdl:4041:8  */
  assign bitheapresult_bh85 = tmp_bitheapresult_bh85_17; // (signal)
  /* fppow16.vhdl:4043:8  */
  assign outres = bitheapresult_bh85; // (signal)
  /* fppow16.vhdl:4048:4  */
  fixrealkcm_freq500_uid84_t0_freq500_uid87 fixrealkcm_freq500_uid84_table0 (
    .x(fixrealkcm_freq500_uid84_a0),
    .y(fixrealkcm_freq500_uid84_table0_n3087));
  /* fppow16.vhdl:4052:44  */
  assign n3090 = fixrealkcm_freq500_uid84_t0[0]; // extract
  /* fppow16.vhdl:4053:44  */
  assign n3091 = fixrealkcm_freq500_uid84_t0[1]; // extract
  /* fppow16.vhdl:4054:44  */
  assign n3092 = fixrealkcm_freq500_uid84_t0[2]; // extract
  /* fppow16.vhdl:4055:44  */
  assign n3093 = fixrealkcm_freq500_uid84_t0[3]; // extract
  /* fppow16.vhdl:4056:44  */
  assign n3094 = fixrealkcm_freq500_uid84_t0[4]; // extract
  /* fppow16.vhdl:4057:44  */
  assign n3095 = fixrealkcm_freq500_uid84_t0[5]; // extract
  /* fppow16.vhdl:4058:44  */
  assign n3096 = fixrealkcm_freq500_uid84_t0[6]; // extract
  /* fppow16.vhdl:4059:44  */
  assign n3097 = fixrealkcm_freq500_uid84_t0[7]; // extract
  /* fppow16.vhdl:4060:44  */
  assign n3098 = fixrealkcm_freq500_uid84_t0[8]; // extract
  /* fppow16.vhdl:4061:44  */
  assign n3099 = fixrealkcm_freq500_uid84_t0[9]; // extract
  /* fppow16.vhdl:4062:45  */
  assign n3100 = fixrealkcm_freq500_uid84_t0[10]; // extract
  /* fppow16.vhdl:4063:45  */
  assign n3101 = fixrealkcm_freq500_uid84_t0[11]; // extract
  /* fppow16.vhdl:4064:45  */
  assign n3102 = fixrealkcm_freq500_uid84_t0[12]; // extract
  /* fppow16.vhdl:4065:45  */
  assign n3103 = fixrealkcm_freq500_uid84_t0[13]; // extract
  /* fppow16.vhdl:4066:45  */
  assign n3104 = fixrealkcm_freq500_uid84_t0[14]; // extract
  /* fppow16.vhdl:4067:45  */
  assign n3105 = fixrealkcm_freq500_uid84_t0[15]; // extract
  /* fppow16.vhdl:4068:45  */
  assign n3106 = fixrealkcm_freq500_uid84_t0[16]; // extract
  /* fppow16.vhdl:4069:45  */
  assign n3107 = fixrealkcm_freq500_uid84_t0[17]; // extract
  /* fppow16.vhdl:4074:44  */
  assign n3108 = {bh85_w17_0, bh85_w16_0};
  /* fppow16.vhdl:4074:57  */
  assign n3109 = {n3108, bh85_w15_0};
  /* fppow16.vhdl:4074:70  */
  assign n3110 = {n3109, bh85_w14_0};
  /* fppow16.vhdl:4074:83  */
  assign n3111 = {n3110, bh85_w13_0};
  /* fppow16.vhdl:4074:96  */
  assign n3112 = {n3111, bh85_w12_0};
  /* fppow16.vhdl:4074:109  */
  assign n3113 = {n3112, bh85_w11_0};
  /* fppow16.vhdl:4074:122  */
  assign n3114 = {n3113, bh85_w10_0};
  /* fppow16.vhdl:4074:135  */
  assign n3115 = {n3114, bh85_w9_0};
  /* fppow16.vhdl:4074:147  */
  assign n3116 = {n3115, bh85_w8_0};
  /* fppow16.vhdl:4074:159  */
  assign n3117 = {n3116, bh85_w7_0};
  /* fppow16.vhdl:4074:171  */
  assign n3118 = {n3117, bh85_w6_0};
  /* fppow16.vhdl:4074:183  */
  assign n3119 = {n3118, bh85_w5_0};
  /* fppow16.vhdl:4074:195  */
  assign n3120 = {n3119, bh85_w4_0};
  /* fppow16.vhdl:4074:207  */
  assign n3121 = {n3120, bh85_w3_0};
  /* fppow16.vhdl:4074:219  */
  assign n3122 = {n3121, bh85_w2_0};
  /* fppow16.vhdl:4074:231  */
  assign n3123 = {n3122, bh85_w1_0};
  /* fppow16.vhdl:4074:243  */
  assign n3124 = {n3123, bh85_w0_0};
endmodule

module fixrealkcm_freq500_uid72
  (input  clk,
   input  [6:0] x,
   output [4:0] r);
  wire [4:0] fixrealkcm_freq500_uid72_a0;
  wire [8:0] fixrealkcm_freq500_uid72_t0;
  wire [8:0] fixrealkcm_freq500_uid72_t0_copy76;
  wire bh73_w0_0;
  wire bh73_w1_0;
  wire bh73_w2_0;
  wire bh73_w3_0;
  wire bh73_w4_0;
  wire bh73_w5_0;
  wire bh73_w6_0;
  wire bh73_w7_0;
  wire bh73_w8_0;
  wire [1:0] fixrealkcm_freq500_uid72_a1;
  wire [3:0] fixrealkcm_freq500_uid72_t1;
  wire [3:0] fixrealkcm_freq500_uid72_t1_copy79;
  wire bh73_w0_1;
  wire bh73_w1_1;
  wire bh73_w2_1;
  wire bh73_w3_1;
  wire [8:0] bitheapfinaladd_bh73_in0;
  wire [8:0] bitheapfinaladd_bh73_in1;
  wire bitheapfinaladd_bh73_cin;
  wire [8:0] bitheapfinaladd_bh73_out;
  wire [8:0] bitheapresult_bh73;
  wire [8:0] outres;
  wire [4:0] n3046;
  wire [8:0] fixrealkcm_freq500_uid72_table0_n3047;
  wire n3050;
  wire n3051;
  wire n3052;
  wire n3053;
  wire n3054;
  wire n3055;
  wire n3056;
  wire n3057;
  wire n3058;
  wire [1:0] n3059;
  wire [3:0] fixrealkcm_freq500_uid72_table1_n3060;
  wire n3063;
  wire n3064;
  wire n3065;
  wire n3066;
  wire [1:0] n3068;
  wire [2:0] n3069;
  wire [3:0] n3070;
  wire [4:0] n3071;
  wire [5:0] n3072;
  wire [6:0] n3073;
  wire [7:0] n3074;
  wire [8:0] n3075;
  wire [5:0] n3077;
  wire [6:0] n3078;
  wire [7:0] n3079;
  wire [8:0] n3080;
  wire [8:0] bitheapfinaladd_bh73_n3082;
  wire [4:0] n3085;
  assign r = n3085; //(module output)
  /* fppow16.vhdl:3867:8  */
  assign fixrealkcm_freq500_uid72_a0 = n3046; // (signal)
  /* fppow16.vhdl:3869:8  */
  assign fixrealkcm_freq500_uid72_t0 = fixrealkcm_freq500_uid72_t0_copy76; // (signal)
  /* fppow16.vhdl:3871:8  */
  assign fixrealkcm_freq500_uid72_t0_copy76 = fixrealkcm_freq500_uid72_table0_n3047; // (signal)
  /* fppow16.vhdl:3873:8  */
  assign bh73_w0_0 = n3050; // (signal)
  /* fppow16.vhdl:3875:8  */
  assign bh73_w1_0 = n3051; // (signal)
  /* fppow16.vhdl:3877:8  */
  assign bh73_w2_0 = n3052; // (signal)
  /* fppow16.vhdl:3879:8  */
  assign bh73_w3_0 = n3053; // (signal)
  /* fppow16.vhdl:3881:8  */
  assign bh73_w4_0 = n3054; // (signal)
  /* fppow16.vhdl:3883:8  */
  assign bh73_w5_0 = n3055; // (signal)
  /* fppow16.vhdl:3885:8  */
  assign bh73_w6_0 = n3056; // (signal)
  /* fppow16.vhdl:3887:8  */
  assign bh73_w7_0 = n3057; // (signal)
  /* fppow16.vhdl:3947:35  */
  assign bh73_w8_0 = n3058; // (signal)
  /* fppow16.vhdl:3891:8  */
  assign fixrealkcm_freq500_uid72_a1 = n3059; // (signal)
  /* fppow16.vhdl:3893:8  */
  assign fixrealkcm_freq500_uid72_t1 = fixrealkcm_freq500_uid72_t1_copy79; // (signal)
  /* fppow16.vhdl:3895:8  */
  assign fixrealkcm_freq500_uid72_t1_copy79 = fixrealkcm_freq500_uid72_table1_n3060; // (signal)
  /* fppow16.vhdl:3897:8  */
  assign bh73_w0_1 = n3063; // (signal)
  /* fppow16.vhdl:3899:8  */
  assign bh73_w1_1 = n3064; // (signal)
  /* fppow16.vhdl:3901:8  */
  assign bh73_w2_1 = n3065; // (signal)
  /* fppow16.vhdl:3903:8  */
  assign bh73_w3_1 = n3066; // (signal)
  /* fppow16.vhdl:3905:8  */
  assign bitheapfinaladd_bh73_in0 = n3075; // (signal)
  /* fppow16.vhdl:3907:8  */
  assign bitheapfinaladd_bh73_in1 = n3080; // (signal)
  /* fppow16.vhdl:3909:8  */
  assign bitheapfinaladd_bh73_cin = 1'b0; // (signal)
  /* fppow16.vhdl:3911:8  */
  assign bitheapfinaladd_bh73_out = bitheapfinaladd_bh73_n3082; // (signal)
  /* fppow16.vhdl:3913:8  */
  assign bitheapresult_bh73 = bitheapfinaladd_bh73_out; // (signal)
  /* fppow16.vhdl:3915:8  */
  assign outres = bitheapresult_bh73; // (signal)
  /* fppow16.vhdl:3919:36  */
  assign n3046 = x[6:2]; // extract
  /* fppow16.vhdl:3920:4  */
  fixrealkcm_freq500_uid72_t0_freq500_uid75 fixrealkcm_freq500_uid72_table0 (
    .x(fixrealkcm_freq500_uid72_a0),
    .y(fixrealkcm_freq500_uid72_table0_n3047));
  /* fppow16.vhdl:3924:44  */
  assign n3050 = fixrealkcm_freq500_uid72_t0[0]; // extract
  /* fppow16.vhdl:3925:44  */
  assign n3051 = fixrealkcm_freq500_uid72_t0[1]; // extract
  /* fppow16.vhdl:3926:44  */
  assign n3052 = fixrealkcm_freq500_uid72_t0[2]; // extract
  /* fppow16.vhdl:3927:44  */
  assign n3053 = fixrealkcm_freq500_uid72_t0[3]; // extract
  /* fppow16.vhdl:3928:44  */
  assign n3054 = fixrealkcm_freq500_uid72_t0[4]; // extract
  /* fppow16.vhdl:3929:44  */
  assign n3055 = fixrealkcm_freq500_uid72_t0[5]; // extract
  /* fppow16.vhdl:3930:44  */
  assign n3056 = fixrealkcm_freq500_uid72_t0[6]; // extract
  /* fppow16.vhdl:3931:44  */
  assign n3057 = fixrealkcm_freq500_uid72_t0[7]; // extract
  /* fppow16.vhdl:3932:44  */
  assign n3058 = fixrealkcm_freq500_uid72_t0[8]; // extract
  /* fppow16.vhdl:3933:36  */
  assign n3059 = x[1:0]; // extract
  /* fppow16.vhdl:3934:4  */
  fixrealkcm_freq500_uid72_t1_freq500_uid78 fixrealkcm_freq500_uid72_table1 (
    .x(fixrealkcm_freq500_uid72_a1),
    .y(fixrealkcm_freq500_uid72_table1_n3060));
  /* fppow16.vhdl:3938:44  */
  assign n3063 = fixrealkcm_freq500_uid72_t1[0]; // extract
  /* fppow16.vhdl:3939:44  */
  assign n3064 = fixrealkcm_freq500_uid72_t1[1]; // extract
  /* fppow16.vhdl:3940:44  */
  assign n3065 = fixrealkcm_freq500_uid72_t1[2]; // extract
  /* fppow16.vhdl:3941:44  */
  assign n3066 = fixrealkcm_freq500_uid72_t1[3]; // extract
  /* fppow16.vhdl:3947:47  */
  assign n3068 = {bh73_w8_0, bh73_w7_0};
  /* fppow16.vhdl:3947:59  */
  assign n3069 = {n3068, bh73_w6_0};
  /* fppow16.vhdl:3947:71  */
  assign n3070 = {n3069, bh73_w5_0};
  /* fppow16.vhdl:3947:83  */
  assign n3071 = {n3070, bh73_w4_0};
  /* fppow16.vhdl:3947:95  */
  assign n3072 = {n3071, bh73_w3_0};
  /* fppow16.vhdl:3947:107  */
  assign n3073 = {n3072, bh73_w2_0};
  /* fppow16.vhdl:3947:119  */
  assign n3074 = {n3073, bh73_w1_0};
  /* fppow16.vhdl:3947:131  */
  assign n3075 = {n3074, bh73_w0_0};
  /* fppow16.vhdl:3948:60  */
  assign n3077 = {5'b00000, bh73_w3_1};
  /* fppow16.vhdl:3948:72  */
  assign n3078 = {n3077, bh73_w2_1};
  /* fppow16.vhdl:3948:84  */
  assign n3079 = {n3078, bh73_w1_1};
  /* fppow16.vhdl:3948:96  */
  assign n3080 = {n3079, bh73_w0_1};
  /* fppow16.vhdl:3951:4  */
  intadder_9_freq500_uid82 bitheapfinaladd_bh73 (
    .clk(clk),
    .x(bitheapfinaladd_bh73_in0),
    .y(bitheapfinaladd_bh73_in1),
    .cin(bitheapfinaladd_bh73_cin),
    .r(bitheapfinaladd_bh73_n3082));
  /* fppow16.vhdl:3959:15  */
  assign n3085 = outres[8:4]; // extract
endmodule

module fixrealkcm_freq500_uid39_t0_freq500_uid42
  (input  [4:0] x,
   output [25:0] y);
  wire [25:0] y0;
  wire [25:0] y1;
  wire n2948;
  wire n2951;
  wire n2954;
  wire n2957;
  wire n2960;
  wire n2963;
  wire n2966;
  wire n2969;
  wire n2972;
  wire n2975;
  wire n2978;
  wire n2981;
  wire n2984;
  wire n2987;
  wire n2990;
  wire n2993;
  wire n2996;
  wire n2999;
  wire n3002;
  wire n3005;
  wire n3008;
  wire n3011;
  wire n3014;
  wire n3017;
  wire n3020;
  wire n3023;
  wire n3026;
  wire n3029;
  wire n3032;
  wire n3035;
  wire n3038;
  wire n3041;
  wire [31:0] n3043;
  reg [25:0] n3044;
  assign y = y1; //(module output)
  /* fppow16.vhdl:438:8  */
  assign y0 = n3044; // (signal)
  /* fppow16.vhdl:440:8  */
  assign y1 = y0; // (signal)
  /* fppow16.vhdl:444:36  */
  assign n2948 = x == 5'b00000;
  /* fppow16.vhdl:445:36  */
  assign n2951 = x == 5'b00001;
  /* fppow16.vhdl:446:36  */
  assign n2954 = x == 5'b00010;
  /* fppow16.vhdl:447:36  */
  assign n2957 = x == 5'b00011;
  /* fppow16.vhdl:448:36  */
  assign n2960 = x == 5'b00100;
  /* fppow16.vhdl:449:36  */
  assign n2963 = x == 5'b00101;
  /* fppow16.vhdl:450:36  */
  assign n2966 = x == 5'b00110;
  /* fppow16.vhdl:451:36  */
  assign n2969 = x == 5'b00111;
  /* fppow16.vhdl:452:36  */
  assign n2972 = x == 5'b01000;
  /* fppow16.vhdl:453:36  */
  assign n2975 = x == 5'b01001;
  /* fppow16.vhdl:454:36  */
  assign n2978 = x == 5'b01010;
  /* fppow16.vhdl:455:36  */
  assign n2981 = x == 5'b01011;
  /* fppow16.vhdl:456:36  */
  assign n2984 = x == 5'b01100;
  /* fppow16.vhdl:457:36  */
  assign n2987 = x == 5'b01101;
  /* fppow16.vhdl:458:36  */
  assign n2990 = x == 5'b01110;
  /* fppow16.vhdl:459:36  */
  assign n2993 = x == 5'b01111;
  /* fppow16.vhdl:460:36  */
  assign n2996 = x == 5'b10000;
  /* fppow16.vhdl:461:36  */
  assign n2999 = x == 5'b10001;
  /* fppow16.vhdl:462:36  */
  assign n3002 = x == 5'b10010;
  /* fppow16.vhdl:463:36  */
  assign n3005 = x == 5'b10011;
  /* fppow16.vhdl:464:36  */
  assign n3008 = x == 5'b10100;
  /* fppow16.vhdl:465:36  */
  assign n3011 = x == 5'b10101;
  /* fppow16.vhdl:466:36  */
  assign n3014 = x == 5'b10110;
  /* fppow16.vhdl:467:36  */
  assign n3017 = x == 5'b10111;
  /* fppow16.vhdl:468:36  */
  assign n3020 = x == 5'b11000;
  /* fppow16.vhdl:469:36  */
  assign n3023 = x == 5'b11001;
  /* fppow16.vhdl:470:36  */
  assign n3026 = x == 5'b11010;
  /* fppow16.vhdl:471:36  */
  assign n3029 = x == 5'b11011;
  /* fppow16.vhdl:472:36  */
  assign n3032 = x == 5'b11100;
  /* fppow16.vhdl:473:36  */
  assign n3035 = x == 5'b11101;
  /* fppow16.vhdl:474:36  */
  assign n3038 = x == 5'b11110;
  /* fppow16.vhdl:475:36  */
  assign n3041 = x == 5'b11111;
  assign n3043 = {n3041, n3038, n3035, n3032, n3029, n3026, n3023, n3020, n3017, n3014, n3011, n3008, n3005, n3002, n2999, n2996, n2993, n2990, n2987, n2984, n2981, n2978, n2975, n2972, n2969, n2966, n2963, n2960, n2957, n2954, n2951, n2948};
  /* fppow16.vhdl:443:4  */
  always @*
    case (n3043)
      32'b10000000000000000000000000000000: n3044 = 26'b10101011111001101000011101;
      32'b01000000000000000000000000000000: n3044 = 26'b10100110010110101111011010;
      32'b00100000000000000000000000000000: n3044 = 26'b10100000110011110110010111;
      32'b00010000000000000000000000000000: n3044 = 26'b10011011010000111101010100;
      32'b00001000000000000000000000000000: n3044 = 26'b10010101101110000100010001;
      32'b00000100000000000000000000000000: n3044 = 26'b10010000001011001011001110;
      32'b00000010000000000000000000000000: n3044 = 26'b10001010101000010010001011;
      32'b00000001000000000000000000000000: n3044 = 26'b10000101000101011001001000;
      32'b00000000100000000000000000000000: n3044 = 26'b01111111100010100000000101;
      32'b00000000010000000000000000000000: n3044 = 26'b01111001111111100111000010;
      32'b00000000001000000000000000000000: n3044 = 26'b01110100011100101101111111;
      32'b00000000000100000000000000000000: n3044 = 26'b01101110111001110100111100;
      32'b00000000000010000000000000000000: n3044 = 26'b01101001010110111011111001;
      32'b00000000000001000000000000000000: n3044 = 26'b01100011110100000010110110;
      32'b00000000000000100000000000000000: n3044 = 26'b01011110010001001001110011;
      32'b00000000000000010000000000000000: n3044 = 26'b01011000101110010000110000;
      32'b00000000000000001000000000000000: n3044 = 26'b01010011001011010111101101;
      32'b00000000000000000100000000000000: n3044 = 26'b01001101101000011110101010;
      32'b00000000000000000010000000000000: n3044 = 26'b01001000000101100101100111;
      32'b00000000000000000001000000000000: n3044 = 26'b01000010100010101100100100;
      32'b00000000000000000000100000000000: n3044 = 26'b00111100111111110011100001;
      32'b00000000000000000000010000000000: n3044 = 26'b00110111011100111010011110;
      32'b00000000000000000000001000000000: n3044 = 26'b00110001111010000001011011;
      32'b00000000000000000000000100000000: n3044 = 26'b00101100010111001000011000;
      32'b00000000000000000000000010000000: n3044 = 26'b00100110110100001111010101;
      32'b00000000000000000000000001000000: n3044 = 26'b00100001010001010110010010;
      32'b00000000000000000000000000100000: n3044 = 26'b00011011101110011101001111;
      32'b00000000000000000000000000010000: n3044 = 26'b00010110001011100100001100;
      32'b00000000000000000000000000001000: n3044 = 26'b00010000101000101011001001;
      32'b00000000000000000000000000000100: n3044 = 26'b00001011000101110010000110;
      32'b00000000000000000000000000000010: n3044 = 26'b00000101100010111001000011;
      32'b00000000000000000000000000000001: n3044 = 26'b00000000000000000000000000;
      default: n3044 = 26'bX;
    endcase
endmodule

module intadder_17_freq500_uid111
  (input  clk,
   input  [16:0] x,
   input  [16:0] y,
   input  cin,
   output [16:0] r);
  wire [16:0] rtmp;
  wire [16:0] x_d1;
  wire [16:0] y_d1;
  wire cin_d1;
  wire cin_d2;
  wire cin_d3;
  wire cin_d4;
  wire cin_d5;
  wire cin_d6;
  wire cin_d7;
  wire cin_d8;
  wire cin_d9;
  wire cin_d10;
  wire cin_d11;
  wire cin_d12;
  wire cin_d13;
  wire cin_d14;
  wire cin_d15;
  wire cin_d16;
  wire cin_d17;
  wire cin_d18;
  wire [16:0] n2922;
  wire [16:0] n2923;
  wire [16:0] n2924;
  reg [16:0] n2925;
  reg [16:0] n2926;
  reg n2927;
  reg n2928;
  reg n2929;
  reg n2930;
  reg n2931;
  reg n2932;
  reg n2933;
  reg n2934;
  reg n2935;
  reg n2936;
  reg n2937;
  reg n2938;
  reg n2939;
  reg n2940;
  reg n2941;
  reg n2942;
  reg n2943;
  reg n2944;
  assign r = rtmp; //(module output)
  /* fppow16.vhdl:4576:8  */
  assign rtmp = n2924; // (signal)
  /* fppow16.vhdl:4578:8  */
  assign x_d1 = n2925; // (signal)
  /* fppow16.vhdl:4580:8  */
  assign y_d1 = n2926; // (signal)
  /* fppow16.vhdl:4582:8  */
  assign cin_d1 = n2927; // (signal)
  /* fppow16.vhdl:4582:16  */
  assign cin_d2 = n2928; // (signal)
  /* fppow16.vhdl:4582:24  */
  assign cin_d3 = n2929; // (signal)
  /* fppow16.vhdl:4582:32  */
  assign cin_d4 = n2930; // (signal)
  /* fppow16.vhdl:4582:40  */
  assign cin_d5 = n2931; // (signal)
  /* fppow16.vhdl:4582:48  */
  assign cin_d6 = n2932; // (signal)
  /* fppow16.vhdl:4582:56  */
  assign cin_d7 = n2933; // (signal)
  /* fppow16.vhdl:4582:64  */
  assign cin_d8 = n2934; // (signal)
  /* fppow16.vhdl:4582:72  */
  assign cin_d9 = n2935; // (signal)
  /* fppow16.vhdl:4582:80  */
  assign cin_d10 = n2936; // (signal)
  /* fppow16.vhdl:4582:89  */
  assign cin_d11 = n2937; // (signal)
  /* fppow16.vhdl:4582:98  */
  assign cin_d12 = n2938; // (signal)
  /* fppow16.vhdl:4582:107  */
  assign cin_d13 = n2939; // (signal)
  /* fppow16.vhdl:4582:116  */
  assign cin_d14 = n2940; // (signal)
  /* fppow16.vhdl:4582:125  */
  assign cin_d15 = n2941; // (signal)
  /* fppow16.vhdl:4582:134  */
  assign cin_d16 = n2942; // (signal)
  /* fppow16.vhdl:4582:143  */
  assign cin_d17 = n2943; // (signal)
  /* fppow16.vhdl:4582:152  */
  assign cin_d18 = n2944; // (signal)
  /* fppow16.vhdl:4610:17  */
  assign n2922 = x_d1 + y_d1;
  /* fppow16.vhdl:4610:24  */
  assign n2923 = {16'b0, cin_d18};  //  uext
  /* fppow16.vhdl:4610:24  */
  assign n2924 = n2922 + n2923;
  /* fppow16.vhdl:4587:10  */
  always @(posedge clk)
    n2925 <= x;
  /* fppow16.vhdl:4587:10  */
  always @(posedge clk)
    n2926 <= y;
  /* fppow16.vhdl:4587:10  */
  always @(posedge clk)
    n2927 <= cin;
  /* fppow16.vhdl:4587:10  */
  always @(posedge clk)
    n2928 <= cin_d1;
  /* fppow16.vhdl:4587:10  */
  always @(posedge clk)
    n2929 <= cin_d2;
  /* fppow16.vhdl:4587:10  */
  always @(posedge clk)
    n2930 <= cin_d3;
  /* fppow16.vhdl:4587:10  */
  always @(posedge clk)
    n2931 <= cin_d4;
  /* fppow16.vhdl:4587:10  */
  always @(posedge clk)
    n2932 <= cin_d5;
  /* fppow16.vhdl:4587:10  */
  always @(posedge clk)
    n2933 <= cin_d6;
  /* fppow16.vhdl:4587:10  */
  always @(posedge clk)
    n2934 <= cin_d7;
  /* fppow16.vhdl:4587:10  */
  always @(posedge clk)
    n2935 <= cin_d8;
  /* fppow16.vhdl:4587:10  */
  always @(posedge clk)
    n2936 <= cin_d9;
  /* fppow16.vhdl:4587:10  */
  always @(posedge clk)
    n2937 <= cin_d10;
  /* fppow16.vhdl:4587:10  */
  always @(posedge clk)
    n2938 <= cin_d11;
  /* fppow16.vhdl:4587:10  */
  always @(posedge clk)
    n2939 <= cin_d12;
  /* fppow16.vhdl:4587:10  */
  always @(posedge clk)
    n2940 <= cin_d13;
  /* fppow16.vhdl:4587:10  */
  always @(posedge clk)
    n2941 <= cin_d14;
  /* fppow16.vhdl:4587:10  */
  always @(posedge clk)
    n2942 <= cin_d15;
  /* fppow16.vhdl:4587:10  */
  always @(posedge clk)
    n2943 <= cin_d16;
  /* fppow16.vhdl:4587:10  */
  always @(posedge clk)
    n2944 <= cin_d17;
endmodule

module exp_5_10_freq500_uid70
  (input  clk,
   input  [16:0] ufixx_i,
   input  xsign,
   output [13:0] expy,
   output [5:0] k);
  wire [16:0] ufixx;
  wire [6:0] xmulin;
  wire [4:0] absk;
  wire [5:0] minusabsk;
  wire [17:0] absklog2;
  wire [12:0] subop1;
  wire [12:0] subop2;
  wire [12:0] y;
  wire [9:0] a;
  wire [2:0] z;
  wire [13:0] expa;
  wire [13:0] expa_copy95;
  wire [2:0] expzm1_p;
  wire [2:0] expzm1_p_copy98;
  wire [3:0] expzm1;
  wire [3:0] expa_t;
  wire [3:0] exparounded0;
  wire [2:0] exparounded;
  wire [4:0] lowerproduct;
  wire [13:0] extendedlowerproduct;
  wire xsign_d1;
  wire xsign_d2;
  wire xsign_d3;
  wire [6:0] n2841;
  wire [4:0] mulinvlog2_n2842;
  wire [5:0] n2846;
  wire [5:0] n2848;
  wire [5:0] n2849;
  wire [5:0] n2851;
  wire [17:0] mullog2_n2852;
  wire [12:0] n2855;
  wire n2856;
  wire [12:0] n2857;
  wire [12:0] n2858;
  wire [12:0] n2859;
  wire [12:0] n2860;
  wire [12:0] n2861;
  wire [12:0] n2862;
  wire [12:0] n2863;
  localparam n2864 = 1'b1;
  wire [12:0] theyadder_n2865;
  wire [9:0] n2868;
  wire [2:0] n2869;
  wire [13:0] expatable_n2870;
  wire [2:0] expzm1table_n2873;
  wire [3:0] n2877;
  wire [3:0] n2878;
  localparam [3:0] n2879 = 4'b0000;
  localparam n2880 = 1'b1;
  wire [3:0] adder_exparounded0_n2881;
  wire [2:0] n2884;
  wire [4:0] thelowerproduct_n2885;
  wire [13:0] n2889;
  localparam n2890 = 1'b0;
  wire [13:0] thefinaladder_n2891;
  reg n2894;
  reg n2895;
  reg n2896;
  assign expy = thefinaladder_n2891; //(module output)
  assign k = n2849; //(module output)
  /* fppow16.vhdl:4434:8  */
  assign xmulin = n2841; // (signal)
  /* fppow16.vhdl:4436:8  */
  assign absk = mulinvlog2_n2842; // (signal)
  /* fppow16.vhdl:4438:8  */
  assign minusabsk = n2848; // (signal)
  /* fppow16.vhdl:4440:8  */
  assign absklog2 = mullog2_n2852; // (signal)
  /* fppow16.vhdl:4442:8  */
  assign subop1 = n2857; // (signal)
  /* fppow16.vhdl:4444:8  */
  assign subop2 = n2861; // (signal)
  /* fppow16.vhdl:4446:8  */
  assign y = theyadder_n2865; // (signal)
  /* fppow16.vhdl:4448:8  */
  assign a = n2868; // (signal)
  /* fppow16.vhdl:4450:8  */
  assign z = n2869; // (signal)
  /* fppow16.vhdl:4452:8  */
  assign expa = expa_copy95; // (signal)
  /* fppow16.vhdl:4454:8  */
  assign expa_copy95 = expatable_n2870; // (signal)
  /* fppow16.vhdl:4456:8  */
  assign expzm1_p = expzm1_p_copy98; // (signal)
  /* fppow16.vhdl:4458:8  */
  assign expzm1_p_copy98 = expzm1table_n2873; // (signal)
  /* fppow16.vhdl:4460:8  */
  assign expzm1 = n2877; // (signal)
  /* fppow16.vhdl:4462:8  */
  assign expa_t = n2878; // (signal)
  /* fppow16.vhdl:4464:8  */
  assign exparounded0 = adder_exparounded0_n2881; // (signal)
  /* fppow16.vhdl:4466:8  */
  assign exparounded = n2884; // (signal)
  /* fppow16.vhdl:4468:8  */
  assign lowerproduct = thelowerproduct_n2885; // (signal)
  /* fppow16.vhdl:4470:8  */
  assign extendedlowerproduct = n2889; // (signal)
  /* fppow16.vhdl:4472:8  */
  assign xsign_d1 = n2894; // (signal)
  /* fppow16.vhdl:4472:18  */
  assign xsign_d2 = n2895; // (signal)
  /* fppow16.vhdl:4472:28  */
  assign xsign_d3 = n2896; // (signal)
  /* fppow16.vhdl:4488:19  */
  assign n2841 = ufixx[16:10]; // extract
  /* fppow16.vhdl:4489:4  */
  fixrealkcm_freq500_uid72 mulinvlog2 (
    .clk(clk),
    .x(xmulin),
    .r(mulinvlog2_n2842));
  /* fppow16.vhdl:4493:44  */
  assign n2846 = {1'b0, absk};
  /* fppow16.vhdl:4493:37  */
  assign n2848 = 6'b000000 - n2846;
  /* fppow16.vhdl:4494:19  */
  assign n2849 = xsign_d3 ? minusabsk : n2851;
  /* fppow16.vhdl:4494:50  */
  assign n2851 = {1'b0, absk};
  /* fppow16.vhdl:4495:4  */
  fixrealkcm_freq500_uid84 mullog2 (
    .clk(clk),
    .x(absk),
    .r(mullog2_n2852));
  /* fppow16.vhdl:4499:36  */
  assign n2855 = ufixx[12:0]; // extract
  /* fppow16.vhdl:4499:64  */
  assign n2856 = ~xsign_d2;
  /* fppow16.vhdl:4499:51  */
  assign n2857 = n2856 ? n2855 : n2859;
  /* fppow16.vhdl:4499:101  */
  assign n2858 = ufixx[12:0]; // extract
  /* fppow16.vhdl:4499:74  */
  assign n2859 = ~n2858;
  /* fppow16.vhdl:4500:22  */
  assign n2860 = absklog2[12:0]; // extract
  /* fppow16.vhdl:4500:36  */
  assign n2861 = xsign_d3 ? n2860 : n2863;
  /* fppow16.vhdl:4500:72  */
  assign n2862 = absklog2[12:0]; // extract
  /* fppow16.vhdl:4500:59  */
  assign n2863 = ~n2862;
  /* fppow16.vhdl:4501:4  */
  intadder_13_freq500_uid92 theyadder (
    .clk(clk),
    .x(subop1),
    .y(subop2),
    .cin(n2864),
    .r(theyadder_n2865));
  /* fppow16.vhdl:4508:10  */
  assign n2868 = y[12:3]; // extract
  /* fppow16.vhdl:4509:10  */
  assign n2869 = y[2:0]; // extract
  /* fppow16.vhdl:4510:4  */
  fixfunctionbytable_freq500_uid94 expatable (
    .x(a),
    .y(expatable_n2870));
  /* fppow16.vhdl:4514:4  */
  fixfunctionbytable_freq500_uid97 expzm1table (
    .x(z),
    .y(expzm1table_n2873));
  /* fppow16.vhdl:4518:15  */
  assign n2877 = {1'b0, expzm1_p};
  /* fppow16.vhdl:4521:18  */
  assign n2878 = expa[13:10]; // extract
  /* fppow16.vhdl:4522:4  */
  intadder_4_freq500_uid102 adder_exparounded0 (
    .clk(clk),
    .x(expa_t),
    .y(n2879),
    .cin(n2880),
    .r(adder_exparounded0_n2881));
  /* fppow16.vhdl:4528:31  */
  assign n2884 = exparounded0[3:1]; // extract
  /* fppow16.vhdl:4529:4  */
  intmultiplier_3x4_5_freq500_uid104 thelowerproduct (
    .clk(clk),
    .x(exparounded),
    .y(expzm1),
    .r(thelowerproduct_n2885));
  /* fppow16.vhdl:4534:50  */
  assign n2889 = {9'b000000000, lowerproduct};
  /* fppow16.vhdl:4536:4  */
  intadder_14_freq500_uid108 thefinaladder (
    .clk(clk),
    .x(expa),
    .y(extendedlowerproduct),
    .cin(n2890),
    .r(thefinaladder_n2891));
  /* fppow16.vhdl:4481:10  */
  always @(posedge clk)
    n2894 <= xsign;
  /* fppow16.vhdl:4481:10  */
  always @(posedge clk)
    n2895 <= xsign_d1;
  /* fppow16.vhdl:4481:10  */
  always @(posedge clk)
    n2896 <= xsign_d2;
endmodule

module leftshifter19_by_max_16_freq500_uid68
  (input  clk,
   input  [18:0] x,
   input  [4:0] s,
   output [34:0] r);
  wire [4:0] ps;
  wire [4:0] ps_d1;
  wire [18:0] level0;
  wire [18:0] level0_d1;
  wire [19:0] level1;
  wire [21:0] level2;
  wire [25:0] level3;
  wire [25:0] level3_d1;
  wire [33:0] level4;
  wire [49:0] level5;
  wire [19:0] n2799;
  wire n2800;
  wire [19:0] n2801;
  wire [19:0] n2803;
  wire [21:0] n2805;
  wire n2806;
  wire [21:0] n2807;
  wire [21:0] n2809;
  wire [25:0] n2811;
  wire n2812;
  wire [25:0] n2813;
  wire [25:0] n2815;
  wire [33:0] n2817;
  wire n2818;
  wire [33:0] n2819;
  wire [33:0] n2821;
  wire [49:0] n2823;
  wire n2824;
  wire [49:0] n2825;
  wire [49:0] n2827;
  wire [34:0] n2828;
  reg [4:0] n2829;
  reg [18:0] n2830;
  reg [25:0] n2831;
  assign r = n2828; //(module output)
  /* fppow16.vhdl:3719:12  */
  assign ps_d1 = n2829; // (signal)
  /* fppow16.vhdl:3721:16  */
  assign level0_d1 = n2830; // (signal)
  /* fppow16.vhdl:3723:8  */
  assign level1 = n2801; // (signal)
  /* fppow16.vhdl:3725:8  */
  assign level2 = n2807; // (signal)
  /* fppow16.vhdl:3727:8  */
  assign level3 = n2813; // (signal)
  /* fppow16.vhdl:3727:16  */
  assign level3_d1 = n2831; // (signal)
  /* fppow16.vhdl:3729:8  */
  assign level4 = n2819; // (signal)
  /* fppow16.vhdl:3731:8  */
  assign level5 = n2825; // (signal)
  /* fppow16.vhdl:3744:23  */
  assign n2799 = {level0_d1, 1'b0};
  /* fppow16.vhdl:3744:52  */
  assign n2800 = ps[0]; // extract
  /* fppow16.vhdl:3744:45  */
  assign n2801 = n2800 ? n2799 : n2803;
  /* fppow16.vhdl:3744:90  */
  assign n2803 = {1'b0, level0_d1};
  /* fppow16.vhdl:3745:20  */
  assign n2805 = {level1, 2'b00};
  /* fppow16.vhdl:3745:49  */
  assign n2806 = ps[1]; // extract
  /* fppow16.vhdl:3745:42  */
  assign n2807 = n2806 ? n2805 : n2809;
  /* fppow16.vhdl:3745:87  */
  assign n2809 = {2'b00, level1};
  /* fppow16.vhdl:3746:20  */
  assign n2811 = {level2, 4'b0000};
  /* fppow16.vhdl:3746:49  */
  assign n2812 = ps[2]; // extract
  /* fppow16.vhdl:3746:42  */
  assign n2813 = n2812 ? n2811 : n2815;
  /* fppow16.vhdl:3746:87  */
  assign n2815 = {4'b0000, level2};
  /* fppow16.vhdl:3747:23  */
  assign n2817 = {level3_d1, 8'b00000000};
  /* fppow16.vhdl:3747:55  */
  assign n2818 = ps_d1[3]; // extract
  /* fppow16.vhdl:3747:45  */
  assign n2819 = n2818 ? n2817 : n2821;
  /* fppow16.vhdl:3747:93  */
  assign n2821 = {8'b00000000, level3_d1};
  /* fppow16.vhdl:3748:20  */
  assign n2823 = {level4, 16'b0000000000000000};
  /* fppow16.vhdl:3748:53  */
  assign n2824 = ps_d1[4]; // extract
  /* fppow16.vhdl:3748:43  */
  assign n2825 = n2824 ? n2823 : n2827;
  /* fppow16.vhdl:3748:92  */
  assign n2827 = {16'b0000000000000000, level4};
  /* fppow16.vhdl:3749:15  */
  assign n2828 = level5[34:0]; // extract
  /* fppow16.vhdl:3736:10  */
  always @(posedge clk)
    n2829 <= ps;
  /* fppow16.vhdl:3736:10  */
  always @(posedge clk)
    n2830 <= level0;
  /* fppow16.vhdl:3736:10  */
  always @(posedge clk)
    n2831 <= level3;
endmodule

module intadder_25_freq500_uid64
  (input  clk,
   input  [24:0] x,
   input  [24:0] y,
   input  cin,
   output [24:0] r);
  wire [24:0] rtmp;
  wire [24:0] x_d1;
  wire [24:0] y_d1;
  wire [24:0] y_d2;
  wire [24:0] y_d3;
  wire [24:0] y_d4;
  wire [24:0] y_d5;
  wire [24:0] y_d6;
  wire [24:0] y_d7;
  wire [24:0] y_d8;
  wire [24:0] y_d9;
  wire [24:0] y_d10;
  wire [24:0] y_d11;
  wire [24:0] y_d12;
  wire cin_d1;
  wire cin_d2;
  wire cin_d3;
  wire cin_d4;
  wire cin_d5;
  wire cin_d6;
  wire cin_d7;
  wire cin_d8;
  wire cin_d9;
  wire cin_d10;
  wire cin_d11;
  wire cin_d12;
  wire [24:0] n2762;
  wire [24:0] n2763;
  wire [24:0] n2764;
  reg [24:0] n2765;
  reg [24:0] n2766;
  reg [24:0] n2767;
  reg [24:0] n2768;
  reg [24:0] n2769;
  reg [24:0] n2770;
  reg [24:0] n2771;
  reg [24:0] n2772;
  reg [24:0] n2773;
  reg [24:0] n2774;
  reg [24:0] n2775;
  reg [24:0] n2776;
  reg [24:0] n2777;
  reg n2778;
  reg n2779;
  reg n2780;
  reg n2781;
  reg n2782;
  reg n2783;
  reg n2784;
  reg n2785;
  reg n2786;
  reg n2787;
  reg n2788;
  reg n2789;
  assign r = rtmp; //(module output)
  /* fppow16.vhdl:3470:8  */
  assign rtmp = n2764; // (signal)
  /* fppow16.vhdl:3472:8  */
  assign x_d1 = n2765; // (signal)
  /* fppow16.vhdl:3474:8  */
  assign y_d1 = n2766; // (signal)
  /* fppow16.vhdl:3474:14  */
  assign y_d2 = n2767; // (signal)
  /* fppow16.vhdl:3474:20  */
  assign y_d3 = n2768; // (signal)
  /* fppow16.vhdl:3474:26  */
  assign y_d4 = n2769; // (signal)
  /* fppow16.vhdl:3474:32  */
  assign y_d5 = n2770; // (signal)
  /* fppow16.vhdl:3474:38  */
  assign y_d6 = n2771; // (signal)
  /* fppow16.vhdl:3474:44  */
  assign y_d7 = n2772; // (signal)
  /* fppow16.vhdl:3474:50  */
  assign y_d8 = n2773; // (signal)
  /* fppow16.vhdl:3474:56  */
  assign y_d9 = n2774; // (signal)
  /* fppow16.vhdl:3474:62  */
  assign y_d10 = n2775; // (signal)
  /* fppow16.vhdl:3474:69  */
  assign y_d11 = n2776; // (signal)
  /* fppow16.vhdl:3474:76  */
  assign y_d12 = n2777; // (signal)
  /* fppow16.vhdl:3476:8  */
  assign cin_d1 = n2778; // (signal)
  /* fppow16.vhdl:3476:16  */
  assign cin_d2 = n2779; // (signal)
  /* fppow16.vhdl:3476:24  */
  assign cin_d3 = n2780; // (signal)
  /* fppow16.vhdl:3476:32  */
  assign cin_d4 = n2781; // (signal)
  /* fppow16.vhdl:3476:40  */
  assign cin_d5 = n2782; // (signal)
  /* fppow16.vhdl:3476:48  */
  assign cin_d6 = n2783; // (signal)
  /* fppow16.vhdl:3476:56  */
  assign cin_d7 = n2784; // (signal)
  /* fppow16.vhdl:3476:64  */
  assign cin_d8 = n2785; // (signal)
  /* fppow16.vhdl:3476:72  */
  assign cin_d9 = n2786; // (signal)
  /* fppow16.vhdl:3476:80  */
  assign cin_d10 = n2787; // (signal)
  /* fppow16.vhdl:3476:89  */
  assign cin_d11 = n2788; // (signal)
  /* fppow16.vhdl:3476:98  */
  assign cin_d12 = n2789; // (signal)
  /* fppow16.vhdl:3509:17  */
  assign n2762 = x_d1 + y_d12;
  /* fppow16.vhdl:3509:25  */
  assign n2763 = {24'b0, cin_d12};  //  uext
  /* fppow16.vhdl:3509:25  */
  assign n2764 = n2762 + n2763;
  /* fppow16.vhdl:3481:10  */
  always @(posedge clk)
    n2765 <= x;
  /* fppow16.vhdl:3481:10  */
  always @(posedge clk)
    n2766 <= y;
  /* fppow16.vhdl:3481:10  */
  always @(posedge clk)
    n2767 <= y_d1;
  /* fppow16.vhdl:3481:10  */
  always @(posedge clk)
    n2768 <= y_d2;
  /* fppow16.vhdl:3481:10  */
  always @(posedge clk)
    n2769 <= y_d3;
  /* fppow16.vhdl:3481:10  */
  always @(posedge clk)
    n2770 <= y_d4;
  /* fppow16.vhdl:3481:10  */
  always @(posedge clk)
    n2771 <= y_d5;
  /* fppow16.vhdl:3481:10  */
  always @(posedge clk)
    n2772 <= y_d6;
  /* fppow16.vhdl:3481:10  */
  always @(posedge clk)
    n2773 <= y_d7;
  /* fppow16.vhdl:3481:10  */
  always @(posedge clk)
    n2774 <= y_d8;
  /* fppow16.vhdl:3481:10  */
  always @(posedge clk)
    n2775 <= y_d9;
  /* fppow16.vhdl:3481:10  */
  always @(posedge clk)
    n2776 <= y_d10;
  /* fppow16.vhdl:3481:10  */
  always @(posedge clk)
    n2777 <= y_d11;
  /* fppow16.vhdl:3481:10  */
  always @(posedge clk)
    n2778 <= cin;
  /* fppow16.vhdl:3481:10  */
  always @(posedge clk)
    n2779 <= cin_d1;
  /* fppow16.vhdl:3481:10  */
  always @(posedge clk)
    n2780 <= cin_d2;
  /* fppow16.vhdl:3481:10  */
  always @(posedge clk)
    n2781 <= cin_d3;
  /* fppow16.vhdl:3481:10  */
  always @(posedge clk)
    n2782 <= cin_d4;
  /* fppow16.vhdl:3481:10  */
  always @(posedge clk)
    n2783 <= cin_d5;
  /* fppow16.vhdl:3481:10  */
  always @(posedge clk)
    n2784 <= cin_d6;
  /* fppow16.vhdl:3481:10  */
  always @(posedge clk)
    n2785 <= cin_d7;
  /* fppow16.vhdl:3481:10  */
  always @(posedge clk)
    n2786 <= cin_d8;
  /* fppow16.vhdl:3481:10  */
  always @(posedge clk)
    n2787 <= cin_d9;
  /* fppow16.vhdl:3481:10  */
  always @(posedge clk)
    n2788 <= cin_d10;
  /* fppow16.vhdl:3481:10  */
  always @(posedge clk)
    n2789 <= cin_d11;
endmodule

module intmultiplier_18x11_21_freq500_uid60
  (input  clk,
   input  [17:0] x,
   input  [10:0] y,
   output [20:0] r);
  wire [17:0] xx;
  wire [10:0] yy;
  wire [10:0] yy_d1;
  wire [10:0] yy_d2;
  wire [10:0] yy_d3;
  wire [10:0] yy_d4;
  wire [10:0] yy_d5;
  wire [10:0] yy_d6;
  wire [10:0] yy_d7;
  wire [10:0] yy_d8;
  wire [10:0] yy_d9;
  wire [10:0] yy_d10;
  wire [28:0] rr;
  wire [28:0] n2718;
  wire [28:0] n2719;
  wire [28:0] n2720;
  wire [20:0] n2721;
  reg [10:0] n2722;
  reg [10:0] n2723;
  reg [10:0] n2724;
  reg [10:0] n2725;
  reg [10:0] n2726;
  reg [10:0] n2727;
  reg [10:0] n2728;
  reg [10:0] n2729;
  reg [10:0] n2730;
  reg [10:0] n2731;
  assign r = n2721; //(module output)
  /* fppow16.vhdl:3410:12  */
  assign yy_d1 = n2722; // (signal)
  /* fppow16.vhdl:3410:19  */
  assign yy_d2 = n2723; // (signal)
  /* fppow16.vhdl:3410:26  */
  assign yy_d3 = n2724; // (signal)
  /* fppow16.vhdl:3410:33  */
  assign yy_d4 = n2725; // (signal)
  /* fppow16.vhdl:3410:40  */
  assign yy_d5 = n2726; // (signal)
  /* fppow16.vhdl:3410:47  */
  assign yy_d6 = n2727; // (signal)
  /* fppow16.vhdl:3410:54  */
  assign yy_d7 = n2728; // (signal)
  /* fppow16.vhdl:3410:61  */
  assign yy_d8 = n2729; // (signal)
  /* fppow16.vhdl:3410:68  */
  assign yy_d9 = n2730; // (signal)
  /* fppow16.vhdl:3410:75  */
  assign yy_d10 = n2731; // (signal)
  /* fppow16.vhdl:3412:8  */
  assign rr = n2720; // (signal)
  /* fppow16.vhdl:3434:12  */
  assign n2718 = {11'b0, xx};  //  uext
  /* fppow16.vhdl:3434:12  */
  assign n2719 = {18'b0, yy_d10};  //  uext
  /* fppow16.vhdl:3434:12  */
  assign n2720 = n2718 * n2719; // umul
  /* fppow16.vhdl:3435:28  */
  assign n2721 = rr[28:8]; // extract
  /* fppow16.vhdl:3417:10  */
  always @(posedge clk)
    n2722 <= yy;
  /* fppow16.vhdl:3417:10  */
  always @(posedge clk)
    n2723 <= yy_d1;
  /* fppow16.vhdl:3417:10  */
  always @(posedge clk)
    n2724 <= yy_d2;
  /* fppow16.vhdl:3417:10  */
  always @(posedge clk)
    n2725 <= yy_d3;
  /* fppow16.vhdl:3417:10  */
  always @(posedge clk)
    n2726 <= yy_d4;
  /* fppow16.vhdl:3417:10  */
  always @(posedge clk)
    n2727 <= yy_d5;
  /* fppow16.vhdl:3417:10  */
  always @(posedge clk)
    n2728 <= yy_d6;
  /* fppow16.vhdl:3417:10  */
  always @(posedge clk)
    n2729 <= yy_d7;
  /* fppow16.vhdl:3417:10  */
  always @(posedge clk)
    n2730 <= yy_d8;
  /* fppow16.vhdl:3417:10  */
  always @(posedge clk)
    n2731 <= yy_d9;
endmodule

module intadder_22_freq500_uid55
  (input  clk,
   input  [21:0] x,
   input  [21:0] y,
   input  cin,
   output [21:0] r);
  wire [21:0] rtmp;
  wire [21:0] x_d1;
  wire [21:0] y_d1;
  wire cin_d1;
  wire cin_d2;
  wire cin_d3;
  wire cin_d4;
  wire cin_d5;
  wire cin_d6;
  wire cin_d7;
  wire cin_d8;
  wire cin_d9;
  wire cin_d10;
  wire [21:0] n2688;
  wire [21:0] n2689;
  wire [21:0] n2690;
  reg [21:0] n2691;
  reg [21:0] n2692;
  reg n2693;
  reg n2694;
  reg n2695;
  reg n2696;
  reg n2697;
  reg n2698;
  reg n2699;
  reg n2700;
  reg n2701;
  reg n2702;
  assign r = rtmp; //(module output)
  /* fppow16.vhdl:2795:8  */
  assign rtmp = n2690; // (signal)
  /* fppow16.vhdl:2797:8  */
  assign x_d1 = n2691; // (signal)
  /* fppow16.vhdl:2799:8  */
  assign y_d1 = n2692; // (signal)
  /* fppow16.vhdl:2801:8  */
  assign cin_d1 = n2693; // (signal)
  /* fppow16.vhdl:2801:16  */
  assign cin_d2 = n2694; // (signal)
  /* fppow16.vhdl:2801:24  */
  assign cin_d3 = n2695; // (signal)
  /* fppow16.vhdl:2801:32  */
  assign cin_d4 = n2696; // (signal)
  /* fppow16.vhdl:2801:40  */
  assign cin_d5 = n2697; // (signal)
  /* fppow16.vhdl:2801:48  */
  assign cin_d6 = n2698; // (signal)
  /* fppow16.vhdl:2801:56  */
  assign cin_d7 = n2699; // (signal)
  /* fppow16.vhdl:2801:64  */
  assign cin_d8 = n2700; // (signal)
  /* fppow16.vhdl:2801:72  */
  assign cin_d9 = n2701; // (signal)
  /* fppow16.vhdl:2801:80  */
  assign cin_d10 = n2702; // (signal)
  /* fppow16.vhdl:2821:17  */
  assign n2688 = x_d1 + y_d1;
  /* fppow16.vhdl:2821:24  */
  assign n2689 = {21'b0, cin_d10};  //  uext
  /* fppow16.vhdl:2821:24  */
  assign n2690 = n2688 + n2689;
  /* fppow16.vhdl:2806:10  */
  always @(posedge clk)
    n2691 <= x;
  /* fppow16.vhdl:2806:10  */
  always @(posedge clk)
    n2692 <= y;
  /* fppow16.vhdl:2806:10  */
  always @(posedge clk)
    n2693 <= cin;
  /* fppow16.vhdl:2806:10  */
  always @(posedge clk)
    n2694 <= cin_d1;
  /* fppow16.vhdl:2806:10  */
  always @(posedge clk)
    n2695 <= cin_d2;
  /* fppow16.vhdl:2806:10  */
  always @(posedge clk)
    n2696 <= cin_d3;
  /* fppow16.vhdl:2806:10  */
  always @(posedge clk)
    n2697 <= cin_d4;
  /* fppow16.vhdl:2806:10  */
  always @(posedge clk)
    n2698 <= cin_d5;
  /* fppow16.vhdl:2806:10  */
  always @(posedge clk)
    n2699 <= cin_d6;
  /* fppow16.vhdl:2806:10  */
  always @(posedge clk)
    n2700 <= cin_d7;
  /* fppow16.vhdl:2806:10  */
  always @(posedge clk)
    n2701 <= cin_d8;
  /* fppow16.vhdl:2806:10  */
  always @(posedge clk)
    n2702 <= cin_d9;
endmodule

module intadder_23_freq500_uid52
  (input  clk,
   input  [22:0] x,
   input  [22:0] y,
   input  cin,
   output [22:0] r);
  wire [22:0] rtmp;
  wire [22:0] x_d1;
  wire [22:0] x_d2;
  wire cin_d1;
  wire cin_d2;
  wire cin_d3;
  wire cin_d4;
  wire cin_d5;
  wire cin_d6;
  wire [22:0] n2660;
  wire [22:0] n2661;
  wire [22:0] n2662;
  reg [22:0] n2663;
  reg [22:0] n2664;
  reg n2665;
  reg n2666;
  reg n2667;
  reg n2668;
  reg n2669;
  reg n2670;
  assign r = rtmp; //(module output)
  /* fppow16.vhdl:2739:8  */
  assign rtmp = n2662; // (signal)
  /* fppow16.vhdl:2741:8  */
  assign x_d1 = n2663; // (signal)
  /* fppow16.vhdl:2741:14  */
  assign x_d2 = n2664; // (signal)
  /* fppow16.vhdl:2743:8  */
  assign cin_d1 = n2665; // (signal)
  /* fppow16.vhdl:2743:16  */
  assign cin_d2 = n2666; // (signal)
  /* fppow16.vhdl:2743:24  */
  assign cin_d3 = n2667; // (signal)
  /* fppow16.vhdl:2743:32  */
  assign cin_d4 = n2668; // (signal)
  /* fppow16.vhdl:2743:40  */
  assign cin_d5 = n2669; // (signal)
  /* fppow16.vhdl:2743:48  */
  assign cin_d6 = n2670; // (signal)
  /* fppow16.vhdl:2759:17  */
  assign n2660 = x_d2 + y;
  /* fppow16.vhdl:2759:21  */
  assign n2661 = {22'b0, cin_d6};  //  uext
  /* fppow16.vhdl:2759:21  */
  assign n2662 = n2660 + n2661;
  /* fppow16.vhdl:2748:10  */
  always @(posedge clk)
    n2663 <= x;
  /* fppow16.vhdl:2748:10  */
  always @(posedge clk)
    n2664 <= x_d1;
  /* fppow16.vhdl:2748:10  */
  always @(posedge clk)
    n2665 <= cin;
  /* fppow16.vhdl:2748:10  */
  always @(posedge clk)
    n2666 <= cin_d1;
  /* fppow16.vhdl:2748:10  */
  always @(posedge clk)
    n2667 <= cin_d2;
  /* fppow16.vhdl:2748:10  */
  always @(posedge clk)
    n2668 <= cin_d3;
  /* fppow16.vhdl:2748:10  */
  always @(posedge clk)
    n2669 <= cin_d4;
  /* fppow16.vhdl:2748:10  */
  always @(posedge clk)
    n2670 <= cin_d5;
endmodule

module rightshifter14_by_max_13_freq500_uid50
  (input  clk,
   input  [13:0] x,
   input  [3:0] s,
   output [26:0] r);
  wire [3:0] ps;
  wire [3:0] ps_d1;
  wire [3:0] ps_d2;
  wire [3:0] ps_d3;
  wire [13:0] level0;
  wire [14:0] level1;
  wire [16:0] level2;
  wire [20:0] level3;
  wire [20:0] level3_d1;
  wire [28:0] level4;
  wire [14:0] n2619;
  wire n2620;
  wire [14:0] n2621;
  wire [14:0] n2623;
  wire [16:0] n2625;
  wire n2626;
  wire [16:0] n2627;
  wire [16:0] n2629;
  wire [20:0] n2631;
  wire n2632;
  wire [20:0] n2633;
  wire [20:0] n2635;
  wire [28:0] n2637;
  wire n2638;
  wire [28:0] n2639;
  wire [28:0] n2641;
  wire [26:0] n2642;
  reg [3:0] n2643;
  reg [3:0] n2644;
  reg [3:0] n2645;
  reg [20:0] n2646;
  assign r = n2642; //(module output)
  /* fppow16.vhdl:2676:12  */
  assign ps_d1 = n2643; // (signal)
  /* fppow16.vhdl:2676:19  */
  assign ps_d2 = n2644; // (signal)
  /* fppow16.vhdl:2676:26  */
  assign ps_d3 = n2645; // (signal)
  /* fppow16.vhdl:2680:8  */
  assign level1 = n2621; // (signal)
  /* fppow16.vhdl:2682:8  */
  assign level2 = n2627; // (signal)
  /* fppow16.vhdl:2684:8  */
  assign level3 = n2633; // (signal)
  /* fppow16.vhdl:2684:16  */
  assign level3_d1 = n2646; // (signal)
  /* fppow16.vhdl:2686:8  */
  assign level4 = n2639; // (signal)
  /* fppow16.vhdl:2700:35  */
  assign n2619 = {1'b0, level0};
  /* fppow16.vhdl:2700:54  */
  assign n2620 = ps_d2[0]; // extract
  /* fppow16.vhdl:2700:44  */
  assign n2621 = n2620 ? n2619 : n2623;
  /* fppow16.vhdl:2700:79  */
  assign n2623 = {level0, 1'b0};
  /* fppow16.vhdl:2701:35  */
  assign n2625 = {2'b00, level1};
  /* fppow16.vhdl:2701:54  */
  assign n2626 = ps_d2[1]; // extract
  /* fppow16.vhdl:2701:44  */
  assign n2627 = n2626 ? n2625 : n2629;
  /* fppow16.vhdl:2701:79  */
  assign n2629 = {level1, 2'b00};
  /* fppow16.vhdl:2702:35  */
  assign n2631 = {4'b0000, level2};
  /* fppow16.vhdl:2702:54  */
  assign n2632 = ps_d2[2]; // extract
  /* fppow16.vhdl:2702:44  */
  assign n2633 = n2632 ? n2631 : n2635;
  /* fppow16.vhdl:2702:79  */
  assign n2635 = {level2, 4'b0000};
  /* fppow16.vhdl:2703:35  */
  assign n2637 = {8'b00000000, level3_d1};
  /* fppow16.vhdl:2703:57  */
  assign n2638 = ps_d3[3]; // extract
  /* fppow16.vhdl:2703:47  */
  assign n2639 = n2638 ? n2637 : n2641;
  /* fppow16.vhdl:2703:85  */
  assign n2641 = {level3_d1, 8'b00000000};
  /* fppow16.vhdl:2704:15  */
  assign n2642 = level4[28:2]; // extract
  /* fppow16.vhdl:2691:10  */
  always @(posedge clk)
    n2643 <= ps;
  /* fppow16.vhdl:2691:10  */
  always @(posedge clk)
    n2644 <= ps_d1;
  /* fppow16.vhdl:2691:10  */
  always @(posedge clk)
    n2645 <= ps_d2;
  /* fppow16.vhdl:2691:10  */
  always @(posedge clk)
    n2646 <= level3;
endmodule

module normalizer_z_35_30_13_freq500_uid48
  (input  clk,
   input  [34:0] x,
   output [3:0] count,
   output [29:0] r);
  wire [34:0] level4;
  wire [34:0] level4_d1;
  wire count3;
  wire count3_d1;
  wire count3_d2;
  wire [34:0] level3;
  wire count2;
  wire count2_d1;
  wire [32:0] level2;
  wire [32:0] level2_d1;
  wire count1;
  wire [30:0] level1;
  wire count0;
  wire [29:0] level0;
  wire [3:0] scount;
  wire [7:0] n2559;
  wire n2561;
  wire n2562;
  wire n2564;
  wire [34:0] n2565;
  wire [26:0] n2566;
  wire [34:0] n2568;
  wire [3:0] n2570;
  wire n2572;
  wire n2573;
  wire [32:0] n2575;
  wire n2576;
  wire [32:0] n2577;
  wire [30:0] n2578;
  wire [32:0] n2580;
  wire [1:0] n2582;
  wire n2584;
  wire n2585;
  wire [30:0] n2587;
  wire n2588;
  wire [30:0] n2589;
  wire [30:0] n2590;
  wire n2592;
  wire n2594;
  wire n2595;
  wire [29:0] n2597;
  wire n2598;
  wire [29:0] n2599;
  wire [29:0] n2600;
  wire [1:0] n2601;
  wire [2:0] n2602;
  wire [3:0] n2603;
  reg [34:0] n2604;
  reg n2605;
  reg n2606;
  reg n2607;
  reg [32:0] n2608;
  assign count = scount; //(module output)
  assign r = level0; //(module output)
  /* fppow16.vhdl:2596:16  */
  assign level4_d1 = n2604; // (signal)
  /* fppow16.vhdl:2598:8  */
  assign count3 = n2562; // (signal)
  /* fppow16.vhdl:2598:16  */
  assign count3_d1 = n2605; // (signal)
  /* fppow16.vhdl:2598:27  */
  assign count3_d2 = n2606; // (signal)
  /* fppow16.vhdl:2600:8  */
  assign level3 = n2565; // (signal)
  /* fppow16.vhdl:2602:8  */
  assign count2 = n2573; // (signal)
  /* fppow16.vhdl:2602:16  */
  assign count2_d1 = n2607; // (signal)
  /* fppow16.vhdl:2604:8  */
  assign level2 = n2577; // (signal)
  /* fppow16.vhdl:2604:16  */
  assign level2_d1 = n2608; // (signal)
  /* fppow16.vhdl:2606:8  */
  assign count1 = n2585; // (signal)
  /* fppow16.vhdl:2608:8  */
  assign level1 = n2589; // (signal)
  /* fppow16.vhdl:2610:8  */
  assign count0 = n2595; // (signal)
  /* fppow16.vhdl:2612:8  */
  assign level0 = n2599; // (signal)
  /* fppow16.vhdl:2614:8  */
  assign scount = n2603; // (signal)
  /* fppow16.vhdl:2628:28  */
  assign n2559 = level4[34:27]; // extract
  /* fppow16.vhdl:2628:43  */
  assign n2561 = n2559 == 8'b00000000;
  /* fppow16.vhdl:2628:17  */
  assign n2562 = n2561 ? 1'b1 : 1'b0;
  /* fppow16.vhdl:2629:50  */
  assign n2564 = ~count3_d1;
  /* fppow16.vhdl:2629:36  */
  assign n2565 = n2564 ? level4_d1 : n2568;
  /* fppow16.vhdl:2629:69  */
  assign n2566 = level4_d1[26:0]; // extract
  /* fppow16.vhdl:2629:83  */
  assign n2568 = {n2566, 8'b00000000};
  /* fppow16.vhdl:2631:28  */
  assign n2570 = level3[34:31]; // extract
  /* fppow16.vhdl:2631:43  */
  assign n2572 = n2570 == 4'b0000;
  /* fppow16.vhdl:2631:17  */
  assign n2573 = n2572 ? 1'b1 : 1'b0;
  /* fppow16.vhdl:2632:19  */
  assign n2575 = level3[34:2]; // extract
  /* fppow16.vhdl:2632:44  */
  assign n2576 = ~count2;
  /* fppow16.vhdl:2632:33  */
  assign n2577 = n2576 ? n2575 : n2580;
  /* fppow16.vhdl:2632:60  */
  assign n2578 = level3[30:0]; // extract
  /* fppow16.vhdl:2632:74  */
  assign n2580 = {n2578, 2'b00};
  /* fppow16.vhdl:2634:31  */
  assign n2582 = level2_d1[32:31]; // extract
  /* fppow16.vhdl:2634:46  */
  assign n2584 = n2582 == 2'b00;
  /* fppow16.vhdl:2634:17  */
  assign n2585 = n2584 ? 1'b1 : 1'b0;
  /* fppow16.vhdl:2635:22  */
  assign n2587 = level2_d1[32:2]; // extract
  /* fppow16.vhdl:2635:47  */
  assign n2588 = ~count1;
  /* fppow16.vhdl:2635:36  */
  assign n2589 = n2588 ? n2587 : n2590;
  /* fppow16.vhdl:2635:66  */
  assign n2590 = level2_d1[30:0]; // extract
  /* fppow16.vhdl:2637:28  */
  assign n2592 = level1[30]; // extract
  /* fppow16.vhdl:2637:43  */
  assign n2594 = n2592 == 1'b0;
  /* fppow16.vhdl:2637:17  */
  assign n2595 = n2594 ? 1'b1 : 1'b0;
  /* fppow16.vhdl:2638:19  */
  assign n2597 = level1[30:1]; // extract
  /* fppow16.vhdl:2638:44  */
  assign n2598 = ~count0;
  /* fppow16.vhdl:2638:33  */
  assign n2599 = n2598 ? n2597 : n2600;
  /* fppow16.vhdl:2638:60  */
  assign n2600 = level1[29:0]; // extract
  /* fppow16.vhdl:2641:24  */
  assign n2601 = {count3_d2, count2_d1};
  /* fppow16.vhdl:2641:36  */
  assign n2602 = {n2601, count1};
  /* fppow16.vhdl:2641:45  */
  assign n2603 = {n2602, count0};
  /* fppow16.vhdl:2619:10  */
  always @(posedge clk)
    n2604 <= level4;
  /* fppow16.vhdl:2619:10  */
  always @(posedge clk)
    n2605 <= count3;
  /* fppow16.vhdl:2619:10  */
  always @(posedge clk)
    n2606 <= count3_d1;
  /* fppow16.vhdl:2619:10  */
  always @(posedge clk)
    n2607 <= count2;
  /* fppow16.vhdl:2619:10  */
  always @(posedge clk)
    n2608 <= level2;
endmodule

module intadder_35_freq500_uid46
  (input  clk,
   input  [34:0] x,
   input  [34:0] y,
   input  cin,
   output [34:0] r);
  wire [34:0] rtmp;
  wire [34:0] x_d1;
  wire [34:0] x_d2;
  wire [34:0] x_d3;
  wire [34:0] x_d4;
  wire [34:0] x_d5;
  wire [34:0] x_d6;
  wire [34:0] y_d1;
  wire cin_d1;
  wire cin_d2;
  wire cin_d3;
  wire cin_d4;
  wire cin_d5;
  wire cin_d6;
  wire cin_d7;
  wire [34:0] n2530;
  wire [34:0] n2531;
  wire [34:0] n2532;
  reg [34:0] n2533;
  reg [34:0] n2534;
  reg [34:0] n2535;
  reg [34:0] n2536;
  reg [34:0] n2537;
  reg [34:0] n2538;
  reg [34:0] n2539;
  reg n2540;
  reg n2541;
  reg n2542;
  reg n2543;
  reg n2544;
  reg n2545;
  reg n2546;
  assign r = rtmp; //(module output)
  /* fppow16.vhdl:2533:8  */
  assign rtmp = n2532; // (signal)
  /* fppow16.vhdl:2535:8  */
  assign x_d1 = n2533; // (signal)
  /* fppow16.vhdl:2535:14  */
  assign x_d2 = n2534; // (signal)
  /* fppow16.vhdl:2535:20  */
  assign x_d3 = n2535; // (signal)
  /* fppow16.vhdl:2535:26  */
  assign x_d4 = n2536; // (signal)
  /* fppow16.vhdl:2535:32  */
  assign x_d5 = n2537; // (signal)
  /* fppow16.vhdl:2535:38  */
  assign x_d6 = n2538; // (signal)
  /* fppow16.vhdl:2537:8  */
  assign y_d1 = n2539; // (signal)
  /* fppow16.vhdl:2539:8  */
  assign cin_d1 = n2540; // (signal)
  /* fppow16.vhdl:2539:16  */
  assign cin_d2 = n2541; // (signal)
  /* fppow16.vhdl:2539:24  */
  assign cin_d3 = n2542; // (signal)
  /* fppow16.vhdl:2539:32  */
  assign cin_d4 = n2543; // (signal)
  /* fppow16.vhdl:2539:40  */
  assign cin_d5 = n2544; // (signal)
  /* fppow16.vhdl:2539:48  */
  assign cin_d6 = n2545; // (signal)
  /* fppow16.vhdl:2539:56  */
  assign cin_d7 = n2546; // (signal)
  /* fppow16.vhdl:2561:17  */
  assign n2530 = x_d6 + y_d1;
  /* fppow16.vhdl:2561:24  */
  assign n2531 = {34'b0, cin_d7};  //  uext
  /* fppow16.vhdl:2561:24  */
  assign n2532 = n2530 + n2531;
  /* fppow16.vhdl:2544:10  */
  always @(posedge clk)
    n2533 <= x;
  /* fppow16.vhdl:2544:10  */
  always @(posedge clk)
    n2534 <= x_d1;
  /* fppow16.vhdl:2544:10  */
  always @(posedge clk)
    n2535 <= x_d2;
  /* fppow16.vhdl:2544:10  */
  always @(posedge clk)
    n2536 <= x_d3;
  /* fppow16.vhdl:2544:10  */
  always @(posedge clk)
    n2537 <= x_d4;
  /* fppow16.vhdl:2544:10  */
  always @(posedge clk)
    n2538 <= x_d5;
  /* fppow16.vhdl:2544:10  */
  always @(posedge clk)
    n2539 <= y;
  /* fppow16.vhdl:2544:10  */
  always @(posedge clk)
    n2540 <= cin;
  /* fppow16.vhdl:2544:10  */
  always @(posedge clk)
    n2541 <= cin_d1;
  /* fppow16.vhdl:2544:10  */
  always @(posedge clk)
    n2542 <= cin_d2;
  /* fppow16.vhdl:2544:10  */
  always @(posedge clk)
    n2543 <= cin_d3;
  /* fppow16.vhdl:2544:10  */
  always @(posedge clk)
    n2544 <= cin_d4;
  /* fppow16.vhdl:2544:10  */
  always @(posedge clk)
    n2545 <= cin_d5;
  /* fppow16.vhdl:2544:10  */
  always @(posedge clk)
    n2546 <= cin_d6;
endmodule

module fixrealkcm_freq500_uid39
  (input  clk,
   input  [4:0] x,
   output [25:0] r);
  wire [4:0] fixrealkcm_freq500_uid39_a0;
  wire [25:0] fixrealkcm_freq500_uid39_t0;
  wire [25:0] fixrealkcm_freq500_uid39_t0_copy43;
  wire [25:0] fixrealkcm_freq500_uid39_t0_copy43_d1;
  wire bh40_w0_0;
  wire bh40_w1_0;
  wire bh40_w2_0;
  wire bh40_w3_0;
  wire bh40_w4_0;
  wire bh40_w5_0;
  wire bh40_w6_0;
  wire bh40_w7_0;
  wire bh40_w8_0;
  wire bh40_w9_0;
  wire bh40_w10_0;
  wire bh40_w11_0;
  wire bh40_w12_0;
  wire bh40_w13_0;
  wire bh40_w14_0;
  wire bh40_w15_0;
  wire bh40_w16_0;
  wire bh40_w17_0;
  wire bh40_w18_0;
  wire bh40_w19_0;
  wire bh40_w20_0;
  wire bh40_w21_0;
  wire bh40_w22_0;
  wire bh40_w23_0;
  wire bh40_w24_0;
  wire bh40_w25_0;
  wire [25:0] tmp_bitheapresult_bh40_25;
  wire [25:0] bitheapresult_bh40;
  wire [25:0] outres;
  wire [25:0] fixrealkcm_freq500_uid39_table0_n2456;
  wire n2459;
  wire n2460;
  wire n2461;
  wire n2462;
  wire n2463;
  wire n2464;
  wire n2465;
  wire n2466;
  wire n2467;
  wire n2468;
  wire n2469;
  wire n2470;
  wire n2471;
  wire n2472;
  wire n2473;
  wire n2474;
  wire n2475;
  wire n2476;
  wire n2477;
  wire n2478;
  wire n2479;
  wire n2480;
  wire n2481;
  wire n2482;
  wire n2483;
  wire n2484;
  wire [1:0] n2485;
  wire [2:0] n2486;
  wire [3:0] n2487;
  wire [4:0] n2488;
  wire [5:0] n2489;
  wire [6:0] n2490;
  wire [7:0] n2491;
  wire [8:0] n2492;
  wire [9:0] n2493;
  wire [10:0] n2494;
  wire [11:0] n2495;
  wire [12:0] n2496;
  wire [13:0] n2497;
  wire [14:0] n2498;
  wire [15:0] n2499;
  wire [16:0] n2500;
  wire [17:0] n2501;
  wire [18:0] n2502;
  wire [19:0] n2503;
  wire [20:0] n2504;
  wire [21:0] n2505;
  wire [22:0] n2506;
  wire [23:0] n2507;
  wire [24:0] n2508;
  wire [25:0] n2509;
  reg [25:0] n2510;
  assign r = outres; //(module output)
  /* fppow16.vhdl:2390:8  */
  assign fixrealkcm_freq500_uid39_t0 = fixrealkcm_freq500_uid39_t0_copy43_d1; // (signal)
  /* fppow16.vhdl:2392:8  */
  assign fixrealkcm_freq500_uid39_t0_copy43 = fixrealkcm_freq500_uid39_table0_n2456; // (signal)
  /* fppow16.vhdl:2392:44  */
  assign fixrealkcm_freq500_uid39_t0_copy43_d1 = n2510; // (signal)
  /* fppow16.vhdl:2394:8  */
  assign bh40_w0_0 = n2459; // (signal)
  /* fppow16.vhdl:2396:8  */
  assign bh40_w1_0 = n2460; // (signal)
  /* fppow16.vhdl:2398:8  */
  assign bh40_w2_0 = n2461; // (signal)
  /* fppow16.vhdl:2400:8  */
  assign bh40_w3_0 = n2462; // (signal)
  /* fppow16.vhdl:2402:8  */
  assign bh40_w4_0 = n2463; // (signal)
  /* fppow16.vhdl:2404:8  */
  assign bh40_w5_0 = n2464; // (signal)
  /* fppow16.vhdl:2406:8  */
  assign bh40_w6_0 = n2465; // (signal)
  /* fppow16.vhdl:2408:8  */
  assign bh40_w7_0 = n2466; // (signal)
  /* fppow16.vhdl:2410:8  */
  assign bh40_w8_0 = n2467; // (signal)
  /* fppow16.vhdl:2412:8  */
  assign bh40_w9_0 = n2468; // (signal)
  /* fppow16.vhdl:2414:8  */
  assign bh40_w10_0 = n2469; // (signal)
  /* fppow16.vhdl:2416:8  */
  assign bh40_w11_0 = n2470; // (signal)
  /* fppow16.vhdl:2418:8  */
  assign bh40_w12_0 = n2471; // (signal)
  /* fppow16.vhdl:2420:8  */
  assign bh40_w13_0 = n2472; // (signal)
  /* fppow16.vhdl:2422:8  */
  assign bh40_w14_0 = n2473; // (signal)
  /* fppow16.vhdl:2424:8  */
  assign bh40_w15_0 = n2474; // (signal)
  /* fppow16.vhdl:2426:8  */
  assign bh40_w16_0 = n2475; // (signal)
  /* fppow16.vhdl:2428:8  */
  assign bh40_w17_0 = n2476; // (signal)
  /* fppow16.vhdl:2430:8  */
  assign bh40_w18_0 = n2477; // (signal)
  /* fppow16.vhdl:2432:8  */
  assign bh40_w19_0 = n2478; // (signal)
  /* fppow16.vhdl:2434:8  */
  assign bh40_w20_0 = n2479; // (signal)
  /* fppow16.vhdl:2436:8  */
  assign bh40_w21_0 = n2480; // (signal)
  /* fppow16.vhdl:2438:8  */
  assign bh40_w22_0 = n2481; // (signal)
  /* fppow16.vhdl:2440:8  */
  assign bh40_w23_0 = n2482; // (signal)
  /* fppow16.vhdl:2442:8  */
  assign bh40_w24_0 = n2483; // (signal)
  /* fppow16.vhdl:2444:8  */
  assign bh40_w25_0 = n2484; // (signal)
  /* fppow16.vhdl:2446:8  */
  assign tmp_bitheapresult_bh40_25 = n2509; // (signal)
  /* fppow16.vhdl:2448:8  */
  assign bitheapresult_bh40 = tmp_bitheapresult_bh40_25; // (signal)
  /* fppow16.vhdl:2450:8  */
  assign outres = bitheapresult_bh40; // (signal)
  /* fppow16.vhdl:2461:4  */
  fixrealkcm_freq500_uid39_t0_freq500_uid42 fixrealkcm_freq500_uid39_table0 (
    .x(fixrealkcm_freq500_uid39_a0),
    .y(fixrealkcm_freq500_uid39_table0_n2456));
  /* fppow16.vhdl:2465:44  */
  assign n2459 = fixrealkcm_freq500_uid39_t0[0]; // extract
  /* fppow16.vhdl:2466:44  */
  assign n2460 = fixrealkcm_freq500_uid39_t0[1]; // extract
  /* fppow16.vhdl:2467:44  */
  assign n2461 = fixrealkcm_freq500_uid39_t0[2]; // extract
  /* fppow16.vhdl:2468:44  */
  assign n2462 = fixrealkcm_freq500_uid39_t0[3]; // extract
  /* fppow16.vhdl:2469:44  */
  assign n2463 = fixrealkcm_freq500_uid39_t0[4]; // extract
  /* fppow16.vhdl:2470:44  */
  assign n2464 = fixrealkcm_freq500_uid39_t0[5]; // extract
  /* fppow16.vhdl:2471:44  */
  assign n2465 = fixrealkcm_freq500_uid39_t0[6]; // extract
  /* fppow16.vhdl:2472:44  */
  assign n2466 = fixrealkcm_freq500_uid39_t0[7]; // extract
  /* fppow16.vhdl:2473:44  */
  assign n2467 = fixrealkcm_freq500_uid39_t0[8]; // extract
  /* fppow16.vhdl:2474:44  */
  assign n2468 = fixrealkcm_freq500_uid39_t0[9]; // extract
  /* fppow16.vhdl:2475:45  */
  assign n2469 = fixrealkcm_freq500_uid39_t0[10]; // extract
  /* fppow16.vhdl:2476:45  */
  assign n2470 = fixrealkcm_freq500_uid39_t0[11]; // extract
  /* fppow16.vhdl:2477:45  */
  assign n2471 = fixrealkcm_freq500_uid39_t0[12]; // extract
  /* fppow16.vhdl:2478:45  */
  assign n2472 = fixrealkcm_freq500_uid39_t0[13]; // extract
  /* fppow16.vhdl:2479:45  */
  assign n2473 = fixrealkcm_freq500_uid39_t0[14]; // extract
  /* fppow16.vhdl:2480:45  */
  assign n2474 = fixrealkcm_freq500_uid39_t0[15]; // extract
  /* fppow16.vhdl:2481:45  */
  assign n2475 = fixrealkcm_freq500_uid39_t0[16]; // extract
  /* fppow16.vhdl:2482:45  */
  assign n2476 = fixrealkcm_freq500_uid39_t0[17]; // extract
  /* fppow16.vhdl:2483:45  */
  assign n2477 = fixrealkcm_freq500_uid39_t0[18]; // extract
  /* fppow16.vhdl:2484:45  */
  assign n2478 = fixrealkcm_freq500_uid39_t0[19]; // extract
  /* fppow16.vhdl:2485:45  */
  assign n2479 = fixrealkcm_freq500_uid39_t0[20]; // extract
  /* fppow16.vhdl:2486:45  */
  assign n2480 = fixrealkcm_freq500_uid39_t0[21]; // extract
  /* fppow16.vhdl:2487:45  */
  assign n2481 = fixrealkcm_freq500_uid39_t0[22]; // extract
  /* fppow16.vhdl:2488:45  */
  assign n2482 = fixrealkcm_freq500_uid39_t0[23]; // extract
  /* fppow16.vhdl:2489:45  */
  assign n2483 = fixrealkcm_freq500_uid39_t0[24]; // extract
  /* fppow16.vhdl:2490:45  */
  assign n2484 = fixrealkcm_freq500_uid39_t0[25]; // extract
  /* fppow16.vhdl:2495:44  */
  assign n2485 = {bh40_w25_0, bh40_w24_0};
  /* fppow16.vhdl:2495:57  */
  assign n2486 = {n2485, bh40_w23_0};
  /* fppow16.vhdl:2495:70  */
  assign n2487 = {n2486, bh40_w22_0};
  /* fppow16.vhdl:2495:83  */
  assign n2488 = {n2487, bh40_w21_0};
  /* fppow16.vhdl:2495:96  */
  assign n2489 = {n2488, bh40_w20_0};
  /* fppow16.vhdl:2495:109  */
  assign n2490 = {n2489, bh40_w19_0};
  /* fppow16.vhdl:2495:122  */
  assign n2491 = {n2490, bh40_w18_0};
  /* fppow16.vhdl:2495:135  */
  assign n2492 = {n2491, bh40_w17_0};
  /* fppow16.vhdl:2495:148  */
  assign n2493 = {n2492, bh40_w16_0};
  /* fppow16.vhdl:2495:161  */
  assign n2494 = {n2493, bh40_w15_0};
  /* fppow16.vhdl:2495:174  */
  assign n2495 = {n2494, bh40_w14_0};
  /* fppow16.vhdl:2495:187  */
  assign n2496 = {n2495, bh40_w13_0};
  /* fppow16.vhdl:2495:200  */
  assign n2497 = {n2496, bh40_w12_0};
  /* fppow16.vhdl:2495:213  */
  assign n2498 = {n2497, bh40_w11_0};
  /* fppow16.vhdl:2495:226  */
  assign n2499 = {n2498, bh40_w10_0};
  /* fppow16.vhdl:2495:239  */
  assign n2500 = {n2499, bh40_w9_0};
  /* fppow16.vhdl:2495:251  */
  assign n2501 = {n2500, bh40_w8_0};
  /* fppow16.vhdl:2495:263  */
  assign n2502 = {n2501, bh40_w7_0};
  /* fppow16.vhdl:2495:275  */
  assign n2503 = {n2502, bh40_w6_0};
  /* fppow16.vhdl:2495:287  */
  assign n2504 = {n2503, bh40_w5_0};
  /* fppow16.vhdl:2495:299  */
  assign n2505 = {n2504, bh40_w4_0};
  /* fppow16.vhdl:2495:311  */
  assign n2506 = {n2505, bh40_w3_0};
  /* fppow16.vhdl:2495:323  */
  assign n2507 = {n2506, bh40_w2_0};
  /* fppow16.vhdl:2495:335  */
  assign n2508 = {n2507, bh40_w1_0};
  /* fppow16.vhdl:2495:347  */
  assign n2509 = {n2508, bh40_w0_0};
  /* fppow16.vhdl:2455:10  */
  always @(posedge clk)
    n2510 <= fixrealkcm_freq500_uid39_t0_copy43;
endmodule

module intadder_30_freq500_uid37
  (input  clk,
   input  [29:0] x,
   input  [29:0] y,
   input  cin,
   output [29:0] r);
  wire [29:0] rtmp;
  wire [29:0] x_d1;
  wire [29:0] x_d2;
  wire [29:0] x_d3;
  wire [29:0] x_d4;
  wire cin_d1;
  wire cin_d2;
  wire cin_d3;
  wire cin_d4;
  wire cin_d5;
  wire cin_d6;
  wire [29:0] n2437;
  wire [29:0] n2438;
  wire [29:0] n2439;
  reg [29:0] n2440;
  reg [29:0] n2441;
  reg [29:0] n2442;
  reg [29:0] n2443;
  reg n2444;
  reg n2445;
  reg n2446;
  reg n2447;
  reg n2448;
  reg n2449;
  assign r = rtmp; //(module output)
  /* fppow16.vhdl:2327:8  */
  assign rtmp = n2439; // (signal)
  /* fppow16.vhdl:2329:8  */
  assign x_d1 = n2440; // (signal)
  /* fppow16.vhdl:2329:14  */
  assign x_d2 = n2441; // (signal)
  /* fppow16.vhdl:2329:20  */
  assign x_d3 = n2442; // (signal)
  /* fppow16.vhdl:2329:26  */
  assign x_d4 = n2443; // (signal)
  /* fppow16.vhdl:2331:8  */
  assign cin_d1 = n2444; // (signal)
  /* fppow16.vhdl:2331:16  */
  assign cin_d2 = n2445; // (signal)
  /* fppow16.vhdl:2331:24  */
  assign cin_d3 = n2446; // (signal)
  /* fppow16.vhdl:2331:32  */
  assign cin_d4 = n2447; // (signal)
  /* fppow16.vhdl:2331:40  */
  assign cin_d5 = n2448; // (signal)
  /* fppow16.vhdl:2331:48  */
  assign cin_d6 = n2449; // (signal)
  /* fppow16.vhdl:2349:17  */
  assign n2437 = x_d4 + y;
  /* fppow16.vhdl:2349:21  */
  assign n2438 = {29'b0, cin_d6};  //  uext
  /* fppow16.vhdl:2349:21  */
  assign n2439 = n2437 + n2438;
  /* fppow16.vhdl:2336:10  */
  always @(posedge clk)
    n2440 <= x;
  /* fppow16.vhdl:2336:10  */
  always @(posedge clk)
    n2441 <= x_d1;
  /* fppow16.vhdl:2336:10  */
  always @(posedge clk)
    n2442 <= x_d2;
  /* fppow16.vhdl:2336:10  */
  always @(posedge clk)
    n2443 <= x_d3;
  /* fppow16.vhdl:2336:10  */
  always @(posedge clk)
    n2444 <= cin;
  /* fppow16.vhdl:2336:10  */
  always @(posedge clk)
    n2445 <= cin_d1;
  /* fppow16.vhdl:2336:10  */
  always @(posedge clk)
    n2446 <= cin_d2;
  /* fppow16.vhdl:2336:10  */
  always @(posedge clk)
    n2447 <= cin_d3;
  /* fppow16.vhdl:2336:10  */
  always @(posedge clk)
    n2448 <= cin_d4;
  /* fppow16.vhdl:2336:10  */
  always @(posedge clk)
    n2449 <= cin_d5;
endmodule

module intadder_30_freq500_uid34
  (input  clk,
   input  [29:0] x,
   input  [29:0] y,
   input  cin,
   output [29:0] r);
  wire cin_1;
  wire cin_1_d1;
  wire cin_1_d2;
  wire [30:0] x_1;
  wire [30:0] x_1_d1;
  wire [30:0] x_1_d2;
  wire [30:0] y_1;
  wire [30:0] y_1_d1;
  wire [30:0] s_1;
  wire [29:0] r_1;
  wire [30:0] n2410;
  wire [30:0] n2412;
  wire [30:0] n2413;
  wire [30:0] n2414;
  wire [30:0] n2415;
  wire [29:0] n2416;
  reg n2417;
  reg n2418;
  reg [30:0] n2419;
  reg [30:0] n2420;
  reg [30:0] n2421;
  assign r = r_1; //(module output)
  /* fppow16.vhdl:2266:15  */
  assign cin_1_d1 = n2417; // (signal)
  /* fppow16.vhdl:2266:25  */
  assign cin_1_d2 = n2418; // (signal)
  /* fppow16.vhdl:2268:8  */
  assign x_1 = n2410; // (signal)
  /* fppow16.vhdl:2268:13  */
  assign x_1_d1 = n2419; // (signal)
  /* fppow16.vhdl:2268:21  */
  assign x_1_d2 = n2420; // (signal)
  /* fppow16.vhdl:2270:8  */
  assign y_1 = n2412; // (signal)
  /* fppow16.vhdl:2270:13  */
  assign y_1_d1 = n2421; // (signal)
  /* fppow16.vhdl:2272:8  */
  assign s_1 = n2415; // (signal)
  /* fppow16.vhdl:2274:8  */
  assign r_1 = n2416; // (signal)
  /* fppow16.vhdl:2288:15  */
  assign n2410 = {1'b0, x};
  /* fppow16.vhdl:2289:15  */
  assign n2412 = {1'b0, y};
  /* fppow16.vhdl:2290:18  */
  assign n2413 = x_1_d2 + y_1_d1;
  /* fppow16.vhdl:2290:27  */
  assign n2414 = {30'b0, cin_1_d2};  //  uext
  /* fppow16.vhdl:2290:27  */
  assign n2415 = n2413 + n2414;
  /* fppow16.vhdl:2291:14  */
  assign n2416 = s_1[29:0]; // extract
  /* fppow16.vhdl:2279:10  */
  always @(posedge clk)
    n2417 <= cin_1;
  /* fppow16.vhdl:2279:10  */
  always @(posedge clk)
    n2418 <= cin_1_d1;
  /* fppow16.vhdl:2279:10  */
  always @(posedge clk)
    n2419 <= x_1;
  /* fppow16.vhdl:2279:10  */
  always @(posedge clk)
    n2420 <= x_1_d1;
  /* fppow16.vhdl:2279:10  */
  always @(posedge clk)
    n2421 <= y_1;
endmodule

module logtable1_freq500_uid30
  (input  [4:0] x,
   output [24:0] y);
  wire [24:0] y0;
  wire [24:0] y1;
  wire n2302;
  wire n2305;
  wire n2308;
  wire n2311;
  wire n2314;
  wire n2317;
  wire n2320;
  wire n2323;
  wire n2326;
  wire n2329;
  wire n2332;
  wire n2335;
  wire n2338;
  wire n2341;
  wire n2344;
  wire n2347;
  wire n2350;
  wire n2353;
  wire n2356;
  wire n2359;
  wire n2362;
  wire n2365;
  wire n2368;
  wire n2371;
  wire n2374;
  wire n2377;
  wire n2380;
  wire n2383;
  wire n2386;
  wire n2389;
  wire n2392;
  wire n2395;
  wire [31:0] n2397;
  reg [24:0] n2398;
  assign y = y1; //(module output)
  /* fppow16.vhdl:366:8  */
  assign y0 = n2398; // (signal)
  /* fppow16.vhdl:368:8  */
  assign y1 = y0; // (signal)
  /* fppow16.vhdl:372:35  */
  assign n2302 = x == 5'b00000;
  /* fppow16.vhdl:373:35  */
  assign n2305 = x == 5'b00001;
  /* fppow16.vhdl:374:35  */
  assign n2308 = x == 5'b00010;
  /* fppow16.vhdl:375:35  */
  assign n2311 = x == 5'b00011;
  /* fppow16.vhdl:376:35  */
  assign n2314 = x == 5'b00100;
  /* fppow16.vhdl:377:35  */
  assign n2317 = x == 5'b00101;
  /* fppow16.vhdl:378:35  */
  assign n2320 = x == 5'b00110;
  /* fppow16.vhdl:379:35  */
  assign n2323 = x == 5'b00111;
  /* fppow16.vhdl:380:35  */
  assign n2326 = x == 5'b01000;
  /* fppow16.vhdl:381:35  */
  assign n2329 = x == 5'b01001;
  /* fppow16.vhdl:382:35  */
  assign n2332 = x == 5'b01010;
  /* fppow16.vhdl:383:35  */
  assign n2335 = x == 5'b01011;
  /* fppow16.vhdl:384:35  */
  assign n2338 = x == 5'b01100;
  /* fppow16.vhdl:385:35  */
  assign n2341 = x == 5'b01101;
  /* fppow16.vhdl:386:35  */
  assign n2344 = x == 5'b01110;
  /* fppow16.vhdl:387:35  */
  assign n2347 = x == 5'b01111;
  /* fppow16.vhdl:388:35  */
  assign n2350 = x == 5'b10000;
  /* fppow16.vhdl:389:35  */
  assign n2353 = x == 5'b10001;
  /* fppow16.vhdl:390:35  */
  assign n2356 = x == 5'b10010;
  /* fppow16.vhdl:391:35  */
  assign n2359 = x == 5'b10011;
  /* fppow16.vhdl:392:35  */
  assign n2362 = x == 5'b10100;
  /* fppow16.vhdl:393:35  */
  assign n2365 = x == 5'b10101;
  /* fppow16.vhdl:394:35  */
  assign n2368 = x == 5'b10110;
  /* fppow16.vhdl:395:35  */
  assign n2371 = x == 5'b10111;
  /* fppow16.vhdl:396:35  */
  assign n2374 = x == 5'b11000;
  /* fppow16.vhdl:397:35  */
  assign n2377 = x == 5'b11001;
  /* fppow16.vhdl:398:35  */
  assign n2380 = x == 5'b11010;
  /* fppow16.vhdl:399:35  */
  assign n2383 = x == 5'b11011;
  /* fppow16.vhdl:400:35  */
  assign n2386 = x == 5'b11100;
  /* fppow16.vhdl:401:35  */
  assign n2389 = x == 5'b11101;
  /* fppow16.vhdl:402:35  */
  assign n2392 = x == 5'b11110;
  /* fppow16.vhdl:403:35  */
  assign n2395 = x == 5'b11111;
  assign n2397 = {n2395, n2392, n2389, n2386, n2383, n2380, n2377, n2374, n2371, n2368, n2365, n2362, n2359, n2356, n2353, n2350, n2347, n2344, n2341, n2338, n2335, n2332, n2329, n2326, n2323, n2320, n2317, n2314, n2311, n2308, n2305, n2302};
  /* fppow16.vhdl:371:4  */
  always @*
    case (n2397)
      32'b10000000000000000000000000000000: n2398 = 25'b1111101110010101111110011;
      32'b01000000000000000000000000000000: n2398 = 25'b1111001101011001001110010;
      32'b00100000000000000000000000000000: n2398 = 25'b1110101100011110100101111;
      32'b00010000000000000000000000000000: n2398 = 25'b1110001011100110000100110;
      32'b00001000000000000000000000000000: n2398 = 25'b1101101010101111101010101;
      32'b00000100000000000000000000000000: n2398 = 25'b1101001001111011010111010;
      32'b00000010000000000000000000000000: n2398 = 25'b1100101001001001001010011;
      32'b00000001000000000000000000000000: n2398 = 25'b1100001000011001000011101;
      32'b00000000100000000000000000000000: n2398 = 25'b1011100111101011000011000;
      32'b00000000010000000000000000000000: n2398 = 25'b1011000110111111000111111;
      32'b00000000001000000000000000000000: n2398 = 25'b1010100110010101010010010;
      32'b00000000000100000000000000000000: n2398 = 25'b1010000101101101100001111;
      32'b00000000000010000000000000000000: n2398 = 25'b1001100101000111110110010;
      32'b00000000000001000000000000000000: n2398 = 25'b1001000100100100001111010;
      32'b00000000000000100000000000000000: n2398 = 25'b1000100100000010101100110;
      32'b00000000000000010000000000000000: n2398 = 25'b1000000011100011001110010;
      32'b00000000000000001000000000000000: n2398 = 25'b0111110011010100010000011;
      32'b00000000000000000100000000000000: n2398 = 25'b0111010010110111110111100;
      32'b00000000000000000010000000000000: n2398 = 25'b0110110010011101100010001;
      32'b00000000000000000001000000000000: n2398 = 25'b0110010010000101010000000;
      32'b00000000000000000000100000000000: n2398 = 25'b0101110001101111000000101;
      32'b00000000000000000000010000000000: n2398 = 25'b0101010001011010110100000;
      32'b00000000000000000000001000000000: n2398 = 25'b0100110001001000101001110;
      32'b00000000000000000000000100000000: n2398 = 25'b0100010000111000100001110;
      32'b00000000000000000000000010000000: n2398 = 25'b0011110000101010011011100;
      32'b00000000000000000000000001000000: n2398 = 25'b0011010000011110010111000;
      32'b00000000000000000000000000100000: n2398 = 25'b0010110000010100010011110;
      32'b00000000000000000000000000010000: n2398 = 25'b0010010000001100010001110;
      32'b00000000000000000000000000001000: n2398 = 25'b0001110000000110010000101;
      32'b00000000000000000000000000000100: n2398 = 25'b0001010000000010010000001;
      32'b00000000000000000000000000000010: n2398 = 25'b0000110000000000010000000;
      32'b00000000000000000000000000000001: n2398 = 25'b0000010000000000010000000;
      default: n2398 = 25'bX;
    endcase
endmodule

module logtable0_freq500_uid27
  (input  [6:0] x,
   output [29:0] y);
  wire [29:0] y0;
  wire [29:0] y1;
  wire n1914;
  wire n1917;
  wire n1920;
  wire n1923;
  wire n1926;
  wire n1929;
  wire n1932;
  wire n1935;
  wire n1938;
  wire n1941;
  wire n1944;
  wire n1947;
  wire n1950;
  wire n1953;
  wire n1956;
  wire n1959;
  wire n1962;
  wire n1965;
  wire n1968;
  wire n1971;
  wire n1974;
  wire n1977;
  wire n1980;
  wire n1983;
  wire n1986;
  wire n1989;
  wire n1992;
  wire n1995;
  wire n1998;
  wire n2001;
  wire n2004;
  wire n2007;
  wire n2010;
  wire n2013;
  wire n2016;
  wire n2019;
  wire n2022;
  wire n2025;
  wire n2028;
  wire n2031;
  wire n2034;
  wire n2037;
  wire n2040;
  wire n2043;
  wire n2046;
  wire n2049;
  wire n2052;
  wire n2055;
  wire n2058;
  wire n2061;
  wire n2064;
  wire n2067;
  wire n2070;
  wire n2073;
  wire n2076;
  wire n2079;
  wire n2082;
  wire n2085;
  wire n2088;
  wire n2091;
  wire n2094;
  wire n2097;
  wire n2100;
  wire n2103;
  wire n2106;
  wire n2109;
  wire n2112;
  wire n2115;
  wire n2118;
  wire n2121;
  wire n2124;
  wire n2127;
  wire n2130;
  wire n2133;
  wire n2136;
  wire n2139;
  wire n2142;
  wire n2145;
  wire n2148;
  wire n2151;
  wire n2154;
  wire n2157;
  wire n2160;
  wire n2163;
  wire n2166;
  wire n2169;
  wire n2172;
  wire n2175;
  wire n2178;
  wire n2181;
  wire n2184;
  wire n2187;
  wire n2190;
  wire n2193;
  wire n2196;
  wire n2199;
  wire n2202;
  wire n2205;
  wire n2208;
  wire n2211;
  wire n2214;
  wire n2217;
  wire n2220;
  wire n2223;
  wire n2226;
  wire n2229;
  wire n2232;
  wire n2235;
  wire n2238;
  wire n2241;
  wire n2244;
  wire n2247;
  wire n2250;
  wire n2253;
  wire n2256;
  wire n2259;
  wire n2262;
  wire n2265;
  wire n2268;
  wire n2271;
  wire n2274;
  wire n2277;
  wire n2280;
  wire n2283;
  wire n2286;
  wire n2289;
  wire n2292;
  wire n2295;
  wire [127:0] n2297;
  reg [29:0] n2298;
  assign y = y1; //(module output)
  /* fppow16.vhdl:198:8  */
  assign y0 = n2298; // (signal)
  /* fppow16.vhdl:200:8  */
  assign y1 = y0; // (signal)
  /* fppow16.vhdl:204:40  */
  assign n1914 = x == 7'b0000000;
  /* fppow16.vhdl:205:40  */
  assign n1917 = x == 7'b0000001;
  /* fppow16.vhdl:206:40  */
  assign n1920 = x == 7'b0000010;
  /* fppow16.vhdl:207:40  */
  assign n1923 = x == 7'b0000011;
  /* fppow16.vhdl:208:40  */
  assign n1926 = x == 7'b0000100;
  /* fppow16.vhdl:209:40  */
  assign n1929 = x == 7'b0000101;
  /* fppow16.vhdl:210:40  */
  assign n1932 = x == 7'b0000110;
  /* fppow16.vhdl:211:40  */
  assign n1935 = x == 7'b0000111;
  /* fppow16.vhdl:212:40  */
  assign n1938 = x == 7'b0001000;
  /* fppow16.vhdl:213:40  */
  assign n1941 = x == 7'b0001001;
  /* fppow16.vhdl:214:40  */
  assign n1944 = x == 7'b0001010;
  /* fppow16.vhdl:215:40  */
  assign n1947 = x == 7'b0001011;
  /* fppow16.vhdl:216:40  */
  assign n1950 = x == 7'b0001100;
  /* fppow16.vhdl:217:40  */
  assign n1953 = x == 7'b0001101;
  /* fppow16.vhdl:218:40  */
  assign n1956 = x == 7'b0001110;
  /* fppow16.vhdl:219:40  */
  assign n1959 = x == 7'b0001111;
  /* fppow16.vhdl:220:40  */
  assign n1962 = x == 7'b0010000;
  /* fppow16.vhdl:221:40  */
  assign n1965 = x == 7'b0010001;
  /* fppow16.vhdl:222:40  */
  assign n1968 = x == 7'b0010010;
  /* fppow16.vhdl:223:40  */
  assign n1971 = x == 7'b0010011;
  /* fppow16.vhdl:224:40  */
  assign n1974 = x == 7'b0010100;
  /* fppow16.vhdl:225:40  */
  assign n1977 = x == 7'b0010101;
  /* fppow16.vhdl:226:40  */
  assign n1980 = x == 7'b0010110;
  /* fppow16.vhdl:227:40  */
  assign n1983 = x == 7'b0010111;
  /* fppow16.vhdl:228:40  */
  assign n1986 = x == 7'b0011000;
  /* fppow16.vhdl:229:40  */
  assign n1989 = x == 7'b0011001;
  /* fppow16.vhdl:230:40  */
  assign n1992 = x == 7'b0011010;
  /* fppow16.vhdl:231:40  */
  assign n1995 = x == 7'b0011011;
  /* fppow16.vhdl:232:40  */
  assign n1998 = x == 7'b0011100;
  /* fppow16.vhdl:233:40  */
  assign n2001 = x == 7'b0011101;
  /* fppow16.vhdl:234:40  */
  assign n2004 = x == 7'b0011110;
  /* fppow16.vhdl:235:40  */
  assign n2007 = x == 7'b0011111;
  /* fppow16.vhdl:236:40  */
  assign n2010 = x == 7'b0100000;
  /* fppow16.vhdl:237:40  */
  assign n2013 = x == 7'b0100001;
  /* fppow16.vhdl:238:40  */
  assign n2016 = x == 7'b0100010;
  /* fppow16.vhdl:239:40  */
  assign n2019 = x == 7'b0100011;
  /* fppow16.vhdl:240:40  */
  assign n2022 = x == 7'b0100100;
  /* fppow16.vhdl:241:40  */
  assign n2025 = x == 7'b0100101;
  /* fppow16.vhdl:242:40  */
  assign n2028 = x == 7'b0100110;
  /* fppow16.vhdl:243:40  */
  assign n2031 = x == 7'b0100111;
  /* fppow16.vhdl:244:40  */
  assign n2034 = x == 7'b0101000;
  /* fppow16.vhdl:245:40  */
  assign n2037 = x == 7'b0101001;
  /* fppow16.vhdl:246:40  */
  assign n2040 = x == 7'b0101010;
  /* fppow16.vhdl:247:40  */
  assign n2043 = x == 7'b0101011;
  /* fppow16.vhdl:248:40  */
  assign n2046 = x == 7'b0101100;
  /* fppow16.vhdl:249:40  */
  assign n2049 = x == 7'b0101101;
  /* fppow16.vhdl:250:40  */
  assign n2052 = x == 7'b0101110;
  /* fppow16.vhdl:251:40  */
  assign n2055 = x == 7'b0101111;
  /* fppow16.vhdl:252:40  */
  assign n2058 = x == 7'b0110000;
  /* fppow16.vhdl:253:40  */
  assign n2061 = x == 7'b0110001;
  /* fppow16.vhdl:254:40  */
  assign n2064 = x == 7'b0110010;
  /* fppow16.vhdl:255:40  */
  assign n2067 = x == 7'b0110011;
  /* fppow16.vhdl:256:40  */
  assign n2070 = x == 7'b0110100;
  /* fppow16.vhdl:257:40  */
  assign n2073 = x == 7'b0110101;
  /* fppow16.vhdl:258:40  */
  assign n2076 = x == 7'b0110110;
  /* fppow16.vhdl:259:40  */
  assign n2079 = x == 7'b0110111;
  /* fppow16.vhdl:260:40  */
  assign n2082 = x == 7'b0111000;
  /* fppow16.vhdl:261:40  */
  assign n2085 = x == 7'b0111001;
  /* fppow16.vhdl:262:40  */
  assign n2088 = x == 7'b0111010;
  /* fppow16.vhdl:263:40  */
  assign n2091 = x == 7'b0111011;
  /* fppow16.vhdl:264:40  */
  assign n2094 = x == 7'b0111100;
  /* fppow16.vhdl:265:40  */
  assign n2097 = x == 7'b0111101;
  /* fppow16.vhdl:266:40  */
  assign n2100 = x == 7'b0111110;
  /* fppow16.vhdl:267:40  */
  assign n2103 = x == 7'b0111111;
  /* fppow16.vhdl:268:40  */
  assign n2106 = x == 7'b1000000;
  /* fppow16.vhdl:269:40  */
  assign n2109 = x == 7'b1000001;
  /* fppow16.vhdl:270:40  */
  assign n2112 = x == 7'b1000010;
  /* fppow16.vhdl:271:40  */
  assign n2115 = x == 7'b1000011;
  /* fppow16.vhdl:272:40  */
  assign n2118 = x == 7'b1000100;
  /* fppow16.vhdl:273:40  */
  assign n2121 = x == 7'b1000101;
  /* fppow16.vhdl:274:40  */
  assign n2124 = x == 7'b1000110;
  /* fppow16.vhdl:275:40  */
  assign n2127 = x == 7'b1000111;
  /* fppow16.vhdl:276:40  */
  assign n2130 = x == 7'b1001000;
  /* fppow16.vhdl:277:40  */
  assign n2133 = x == 7'b1001001;
  /* fppow16.vhdl:278:40  */
  assign n2136 = x == 7'b1001010;
  /* fppow16.vhdl:279:40  */
  assign n2139 = x == 7'b1001011;
  /* fppow16.vhdl:280:40  */
  assign n2142 = x == 7'b1001100;
  /* fppow16.vhdl:281:40  */
  assign n2145 = x == 7'b1001101;
  /* fppow16.vhdl:282:40  */
  assign n2148 = x == 7'b1001110;
  /* fppow16.vhdl:283:40  */
  assign n2151 = x == 7'b1001111;
  /* fppow16.vhdl:284:40  */
  assign n2154 = x == 7'b1010000;
  /* fppow16.vhdl:285:40  */
  assign n2157 = x == 7'b1010001;
  /* fppow16.vhdl:286:40  */
  assign n2160 = x == 7'b1010010;
  /* fppow16.vhdl:287:40  */
  assign n2163 = x == 7'b1010011;
  /* fppow16.vhdl:288:40  */
  assign n2166 = x == 7'b1010100;
  /* fppow16.vhdl:289:40  */
  assign n2169 = x == 7'b1010101;
  /* fppow16.vhdl:290:40  */
  assign n2172 = x == 7'b1010110;
  /* fppow16.vhdl:291:40  */
  assign n2175 = x == 7'b1010111;
  /* fppow16.vhdl:292:40  */
  assign n2178 = x == 7'b1011000;
  /* fppow16.vhdl:293:40  */
  assign n2181 = x == 7'b1011001;
  /* fppow16.vhdl:294:40  */
  assign n2184 = x == 7'b1011010;
  /* fppow16.vhdl:295:40  */
  assign n2187 = x == 7'b1011011;
  /* fppow16.vhdl:296:40  */
  assign n2190 = x == 7'b1011100;
  /* fppow16.vhdl:297:40  */
  assign n2193 = x == 7'b1011101;
  /* fppow16.vhdl:298:40  */
  assign n2196 = x == 7'b1011110;
  /* fppow16.vhdl:299:40  */
  assign n2199 = x == 7'b1011111;
  /* fppow16.vhdl:300:40  */
  assign n2202 = x == 7'b1100000;
  /* fppow16.vhdl:301:40  */
  assign n2205 = x == 7'b1100001;
  /* fppow16.vhdl:302:40  */
  assign n2208 = x == 7'b1100010;
  /* fppow16.vhdl:303:40  */
  assign n2211 = x == 7'b1100011;
  /* fppow16.vhdl:304:40  */
  assign n2214 = x == 7'b1100100;
  /* fppow16.vhdl:305:40  */
  assign n2217 = x == 7'b1100101;
  /* fppow16.vhdl:306:40  */
  assign n2220 = x == 7'b1100110;
  /* fppow16.vhdl:307:40  */
  assign n2223 = x == 7'b1100111;
  /* fppow16.vhdl:308:40  */
  assign n2226 = x == 7'b1101000;
  /* fppow16.vhdl:309:40  */
  assign n2229 = x == 7'b1101001;
  /* fppow16.vhdl:310:40  */
  assign n2232 = x == 7'b1101010;
  /* fppow16.vhdl:311:40  */
  assign n2235 = x == 7'b1101011;
  /* fppow16.vhdl:312:40  */
  assign n2238 = x == 7'b1101100;
  /* fppow16.vhdl:313:40  */
  assign n2241 = x == 7'b1101101;
  /* fppow16.vhdl:314:40  */
  assign n2244 = x == 7'b1101110;
  /* fppow16.vhdl:315:40  */
  assign n2247 = x == 7'b1101111;
  /* fppow16.vhdl:316:40  */
  assign n2250 = x == 7'b1110000;
  /* fppow16.vhdl:317:40  */
  assign n2253 = x == 7'b1110001;
  /* fppow16.vhdl:318:40  */
  assign n2256 = x == 7'b1110010;
  /* fppow16.vhdl:319:40  */
  assign n2259 = x == 7'b1110011;
  /* fppow16.vhdl:320:40  */
  assign n2262 = x == 7'b1110100;
  /* fppow16.vhdl:321:40  */
  assign n2265 = x == 7'b1110101;
  /* fppow16.vhdl:322:40  */
  assign n2268 = x == 7'b1110110;
  /* fppow16.vhdl:323:40  */
  assign n2271 = x == 7'b1110111;
  /* fppow16.vhdl:324:40  */
  assign n2274 = x == 7'b1111000;
  /* fppow16.vhdl:325:40  */
  assign n2277 = x == 7'b1111001;
  /* fppow16.vhdl:326:40  */
  assign n2280 = x == 7'b1111010;
  /* fppow16.vhdl:327:40  */
  assign n2283 = x == 7'b1111011;
  /* fppow16.vhdl:328:40  */
  assign n2286 = x == 7'b1111100;
  /* fppow16.vhdl:329:40  */
  assign n2289 = x == 7'b1111101;
  /* fppow16.vhdl:330:40  */
  assign n2292 = x == 7'b1111110;
  /* fppow16.vhdl:331:40  */
  assign n2295 = x == 7'b1111111;
  assign n2297 = {n2295, n2292, n2289, n2286, n2283, n2280, n2277, n2274, n2271, n2268, n2265, n2262, n2259, n2256, n2253, n2250, n2247, n2244, n2241, n2238, n2235, n2232, n2229, n2226, n2223, n2220, n2217, n2214, n2211, n2208, n2205, n2202, n2199, n2196, n2193, n2190, n2187, n2184, n2181, n2178, n2175, n2172, n2169, n2166, n2163, n2160, n2157, n2154, n2151, n2148, n2145, n2142, n2139, n2136, n2133, n2130, n2127, n2124, n2121, n2118, n2115, n2112, n2109, n2106, n2103, n2100, n2097, n2094, n2091, n2088, n2085, n2082, n2079, n2076, n2073, n2070, n2067, n2064, n2061, n2058, n2055, n2052, n2049, n2046, n2043, n2040, n2037, n2034, n2031, n2028, n2025, n2022, n2019, n2016, n2013, n2010, n2007, n2004, n2001, n1998, n1995, n1992, n1989, n1986, n1983, n1980, n1977, n1974, n1971, n1968, n1965, n1962, n1959, n1956, n1953, n1950, n1947, n1944, n1941, n1938, n1935, n1932, n1929, n1926, n1923, n1920, n1917, n1914};
  /* fppow16.vhdl:203:4  */
  always @*
    case (n2297)
      128'b10000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2298 = 30'b111111011100000111111101010110;
      128'b01000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2298 = 30'b111110111100011111101010111010;
      128'b00100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2298 = 30'b111110111100011111101010111010;
      128'b00010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2298 = 30'b111110011101000110111001010000;
      128'b00001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2298 = 30'b111110011101000110111001010000;
      128'b00000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2298 = 30'b111101111101111101011001001111;
      128'b00000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2298 = 30'b111101111101111101011001001111;
      128'b00000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2298 = 30'b111101011111000010111100001001;
      128'b00000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2298 = 30'b111101011111000010111100001001;
      128'b00000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2298 = 30'b111101000000010111010011100001;
      128'b00000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2298 = 30'b111101000000010111010011100001;
      128'b00000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2298 = 30'b111100100001111010010001010010;
      128'b00000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2298 = 30'b111100100001111010010001010010;
      128'b00000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2298 = 30'b111100000011101011100111101000;
      128'b00000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2298 = 30'b111100000011101011100111101000;
      128'b00000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2298 = 30'b111011100101101011001001000100;
      128'b00000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2298 = 30'b111011000111111000101000011010;
      128'b00000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2298 = 30'b111011000111111000101000011010;
      128'b00000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2298 = 30'b111010101010010011111000110000;
      128'b00000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2298 = 30'b111010101010010011111000110000;
      128'b00000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2298 = 30'b111010001100111100101101011101;
      128'b00000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2298 = 30'b111001101111110010111010001010;
      128'b00000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2298 = 30'b111001101111110010111010001010;
      128'b00000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2298 = 30'b111001010010110110010010110001;
      128'b00000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2298 = 30'b111001010010110110010010110001;
      128'b00000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2298 = 30'b111000110110000110101011011100;
      128'b00000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2298 = 30'b111000011001100011111000100100;
      128'b00000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2298 = 30'b111000011001100011111000100100;
      128'b00000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2298 = 30'b110111111101001101101110110100;
      128'b00000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2298 = 30'b110111111101001101101110110100;
      128'b00000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2298 = 30'b110111100001000100000011000010;
      128'b00000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2298 = 30'b110111000101000110101010010110;
      128'b00000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2298 = 30'b110111000101000110101010010110;
      128'b00000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2298 = 30'b110110101001010101011010000100;
      128'b00000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2298 = 30'b110110001101110000000111110000;
      128'b00000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2298 = 30'b110110001101110000000111110000;
      128'b00000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2298 = 30'b110101110010010110101001001010;
      128'b00000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2298 = 30'b110101010111001000110100001110;
      128'b00000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2298 = 30'b110100111100000110011111001000;
      128'b00000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2298 = 30'b110100111100000110011111001000;
      128'b00000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2298 = 30'b110100100001001111100000001100;
      128'b00000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2298 = 30'b110100000110100011101101111111;
      128'b00000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2298 = 30'b110100000110100011101101111111;
      128'b00000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2298 = 30'b110011101100000010111111001110;
      128'b00000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2298 = 30'b110011010001101101001010110010;
      128'b00000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2298 = 30'b110010110111100010000111110000;
      128'b00000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2298 = 30'b110010110111100010000111110000;
      128'b00000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000: n2298 = 30'b110010011101100001101101011001;
      128'b00000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000: n2298 = 30'b110010000011101011110011000110;
      128'b00000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000: n2298 = 30'b110001101010000000010000011100;
      128'b00000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000: n2298 = 30'b110001101010000000010000011100;
      128'b00000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000: n2298 = 30'b110001010000011110111101001010;
      128'b00000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000: n2298 = 30'b110000110111000111110001001001;
      128'b00000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000: n2298 = 30'b110000011101111010100100011010;
      128'b00000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000: n2298 = 30'b110000000100110111001111001001;
      128'b00000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000: n2298 = 30'b110000000100110111001111001001;
      128'b00000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000: n2298 = 30'b101111101011111101101001101100;
      128'b00000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000: n2298 = 30'b101111010011001101101100011110;
      128'b00000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000: n2298 = 30'b101110111010100111010000000110;
      128'b00000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000: n2298 = 30'b101110100010001010001101010100;
      128'b00000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000: n2298 = 30'b101110001001110110011100111110;
      128'b00000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000: n2298 = 30'b101110001001110110011100111110;
      128'b00000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000: n2298 = 30'b101101110001101011111000000100;
      128'b00000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000: n2298 = 30'b101101011001101010010111101100;
      128'b00000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000: n2298 = 30'b011001011000111010001101000011;
      128'b00000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000: n2298 = 30'b011000101001100011100110101000;
      128'b00000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000: n2298 = 30'b011000101001100011100110101000;
      128'b00000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000: n2298 = 30'b010111111010101111101000111100;
      128'b00000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000: n2298 = 30'b010111111010101111101000111100;
      128'b00000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000: n2298 = 30'b010111001100011101100001110111;
      128'b00000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000: n2298 = 30'b010111001100011101100001110111;
      128'b00000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000: n2298 = 30'b010110011110101100100000111110;
      128'b00000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000: n2298 = 30'b010110011110101100100000111110;
      128'b00000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000: n2298 = 30'b010101110001011011110111100000;
      128'b00000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000: n2298 = 30'b010101110001011011110111100000;
      128'b00000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000: n2298 = 30'b010101000100101010111000000111;
      128'b00000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000: n2298 = 30'b010101000100101010111000000111;
      128'b00000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000: n2298 = 30'b010100011000011000110111000010;
      128'b00000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000: n2298 = 30'b010100011000011000110111000010;
      128'b00000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000: n2298 = 30'b010011101100100101001001110111;
      128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000: n2298 = 30'b010011101100100101001001110111;
      128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000: n2298 = 30'b010011000001001111000111100010;
      128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000: n2298 = 30'b010011000001001111000111100010;
      128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000: n2298 = 30'b010010010110010110001000010001;
      128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000: n2298 = 30'b010010010110010110001000010001;
      128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000: n2298 = 30'b010001101011111001100101100100;
      128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000: n2298 = 30'b010001101011111001100101100100;
      128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000: n2298 = 30'b010001000001111000111010000010;
      128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000: n2298 = 30'b010000011000010011100001100000;
      128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000: n2298 = 30'b010000011000010011100001100000;
      128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000: n2298 = 30'b001111101111001000111000110110;
      128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000: n2298 = 30'b001111101111001000111000110110;
      128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000: n2298 = 30'b001111000110011000011110000000;
      128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000: n2298 = 30'b001110011110000001101111111001;
      128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000: n2298 = 30'b001110011110000001101111111001;
      128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000: n2298 = 30'b001101110110000100001110011100;
      128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000: n2298 = 30'b001101001110011111011010011110;
      128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000: n2298 = 30'b001101001110011111011010011110;
      128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000: n2298 = 30'b001100100111010010110101101110;
      128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000: n2298 = 30'b001100000000011110000010110011;
      128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000: n2298 = 30'b001100000000011110000010110011;
      128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000: n2298 = 30'b001011011010000000100101000110;
      128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000: n2298 = 30'b001010110011111010000000110110;
      128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000: n2298 = 30'b001010110011111010000000110110;
      128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000: n2298 = 30'b001010001110001001111011000010;
      128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000: n2298 = 30'b001001101000101111111001011000;
      128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000: n2298 = 30'b001001101000101111111001011000;
      128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000: n2298 = 30'b001001000011101011100010010101;
      128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000: n2298 = 30'b001000011110111100011101000001;
      128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000: n2298 = 30'b000111111010100010010001001110;
      128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000: n2298 = 30'b000111111010100010010001001110;
      128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000: n2298 = 30'b000111010110011100100111011001;
      128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000: n2298 = 30'b000110110010101011001000100011;
      128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000: n2298 = 30'b000110001111001101011110010111;
      128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000: n2298 = 30'b000101101100000011010011000011;
      128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000: n2298 = 30'b000101001001001100010001010111;
      128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000: n2298 = 30'b000101001001001100010001010111;
      128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000: n2298 = 30'b000100100110101000000100101001;
      128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000: n2298 = 30'b000100000100010110011000101101;
      128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000: n2298 = 30'b000011100010010110111001111010;
      128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000: n2298 = 30'b000011000000101001010101000011;
      128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000: n2298 = 30'b000010011111001101010111011010;
      128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000: n2298 = 30'b000001111110000010101110110001;
      128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000: n2298 = 30'b000001011101001001001001010011;
      128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000: n2298 = 30'b000000111100100000010101100110;
      128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100: n2298 = 30'b000000011100001000000010101100;
      128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010: n2298 = 30'b111111111100000000000000000000;
      128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001: n2298 = 30'b111111111100000000000000000000;
      default: n2298 = 30'bX;
    endcase
endmodule

module intadder_21_freq500_uid25
  (input  clk,
   input  [20:0] x,
   input  [20:0] y,
   input  cin,
   output [20:0] r);
  wire [20:0] rtmp;
  wire [20:0] x_d1;
  wire [20:0] x_d2;
  wire [20:0] x_d3;
  wire [20:0] y_d1;
  wire cin_d1;
  wire cin_d2;
  wire cin_d3;
  wire cin_d4;
  wire cin_d5;
  wire cin_d6;
  wire [20:0] n1898;
  wire [20:0] n1899;
  wire [20:0] n1900;
  reg [20:0] n1901;
  reg [20:0] n1902;
  reg [20:0] n1903;
  reg [20:0] n1904;
  reg n1905;
  reg n1906;
  reg n1907;
  reg n1908;
  reg n1909;
  reg n1910;
  assign r = rtmp; //(module output)
  /* fppow16.vhdl:2206:8  */
  assign rtmp = n1900; // (signal)
  /* fppow16.vhdl:2208:8  */
  assign x_d1 = n1901; // (signal)
  /* fppow16.vhdl:2208:14  */
  assign x_d2 = n1902; // (signal)
  /* fppow16.vhdl:2208:20  */
  assign x_d3 = n1903; // (signal)
  /* fppow16.vhdl:2210:8  */
  assign y_d1 = n1904; // (signal)
  /* fppow16.vhdl:2212:8  */
  assign cin_d1 = n1905; // (signal)
  /* fppow16.vhdl:2212:16  */
  assign cin_d2 = n1906; // (signal)
  /* fppow16.vhdl:2212:24  */
  assign cin_d3 = n1907; // (signal)
  /* fppow16.vhdl:2212:32  */
  assign cin_d4 = n1908; // (signal)
  /* fppow16.vhdl:2212:40  */
  assign cin_d5 = n1909; // (signal)
  /* fppow16.vhdl:2212:48  */
  assign cin_d6 = n1910; // (signal)
  /* fppow16.vhdl:2230:17  */
  assign n1898 = x_d3 + y_d1;
  /* fppow16.vhdl:2230:24  */
  assign n1899 = {20'b0, cin_d6};  //  uext
  /* fppow16.vhdl:2230:24  */
  assign n1900 = n1898 + n1899;
  /* fppow16.vhdl:2217:10  */
  always @(posedge clk)
    n1901 <= x;
  /* fppow16.vhdl:2217:10  */
  always @(posedge clk)
    n1902 <= x_d1;
  /* fppow16.vhdl:2217:10  */
  always @(posedge clk)
    n1903 <= x_d2;
  /* fppow16.vhdl:2217:10  */
  always @(posedge clk)
    n1904 <= y;
  /* fppow16.vhdl:2217:10  */
  always @(posedge clk)
    n1905 <= cin;
  /* fppow16.vhdl:2217:10  */
  always @(posedge clk)
    n1906 <= cin_d1;
  /* fppow16.vhdl:2217:10  */
  always @(posedge clk)
    n1907 <= cin_d2;
  /* fppow16.vhdl:2217:10  */
  always @(posedge clk)
    n1908 <= cin_d3;
  /* fppow16.vhdl:2217:10  */
  always @(posedge clk)
    n1909 <= cin_d4;
  /* fppow16.vhdl:2217:10  */
  always @(posedge clk)
    n1910 <= cin_d5;
endmodule

module intadder_21_freq500_uid22
  (input  clk,
   input  [20:0] x,
   input  [20:0] y,
   input  cin,
   output [20:0] r);
  wire cin_1;
  wire cin_1_d1;
  wire cin_1_d2;
  wire cin_1_d3;
  wire [21:0] x_1;
  wire [21:0] x_1_d1;
  wire [21:0] y_1;
  wire [21:0] y_1_d1;
  wire [21:0] s_1;
  wire [20:0] r_1;
  wire [21:0] n1871;
  wire [21:0] n1873;
  wire [21:0] n1874;
  wire [21:0] n1875;
  wire [21:0] n1876;
  wire [20:0] n1877;
  reg n1878;
  reg n1879;
  reg n1880;
  reg [21:0] n1881;
  reg [21:0] n1882;
  assign r = r_1; //(module output)
  /* fppow16.vhdl:2145:15  */
  assign cin_1_d1 = n1878; // (signal)
  /* fppow16.vhdl:2145:25  */
  assign cin_1_d2 = n1879; // (signal)
  /* fppow16.vhdl:2145:35  */
  assign cin_1_d3 = n1880; // (signal)
  /* fppow16.vhdl:2147:8  */
  assign x_1 = n1871; // (signal)
  /* fppow16.vhdl:2147:13  */
  assign x_1_d1 = n1881; // (signal)
  /* fppow16.vhdl:2149:8  */
  assign y_1 = n1873; // (signal)
  /* fppow16.vhdl:2149:13  */
  assign y_1_d1 = n1882; // (signal)
  /* fppow16.vhdl:2151:8  */
  assign s_1 = n1876; // (signal)
  /* fppow16.vhdl:2153:8  */
  assign r_1 = n1877; // (signal)
  /* fppow16.vhdl:2167:15  */
  assign n1871 = {1'b0, x};
  /* fppow16.vhdl:2168:15  */
  assign n1873 = {1'b0, y};
  /* fppow16.vhdl:2169:18  */
  assign n1874 = x_1_d1 + y_1_d1;
  /* fppow16.vhdl:2169:27  */
  assign n1875 = {21'b0, cin_1_d3};  //  uext
  /* fppow16.vhdl:2169:27  */
  assign n1876 = n1874 + n1875;
  /* fppow16.vhdl:2170:14  */
  assign n1877 = s_1[20:0]; // extract
  /* fppow16.vhdl:2158:10  */
  always @(posedge clk)
    n1878 <= cin_1;
  /* fppow16.vhdl:2158:10  */
  always @(posedge clk)
    n1879 <= cin_1_d1;
  /* fppow16.vhdl:2158:10  */
  always @(posedge clk)
    n1880 <= cin_1_d2;
  /* fppow16.vhdl:2158:10  */
  always @(posedge clk)
    n1881 <= x_1;
  /* fppow16.vhdl:2158:10  */
  always @(posedge clk)
    n1882 <= y_1;
endmodule

module intadder_21_freq500_uid19
  (input  clk,
   input  [20:0] x,
   input  [20:0] y,
   input  cin,
   output [20:0] r);
  wire cin_1;
  wire cin_1_d1;
  wire cin_1_d2;
  wire [21:0] x_1;
  wire [21:0] x_1_d1;
  wire [21:0] y_1;
  wire [21:0] y_1_d1;
  wire [21:0] s_1;
  wire [20:0] r_1;
  wire [21:0] n1849;
  wire [21:0] n1851;
  wire [21:0] n1852;
  wire [21:0] n1853;
  wire [21:0] n1854;
  wire [20:0] n1855;
  reg n1856;
  reg n1857;
  reg [21:0] n1858;
  reg [21:0] n1859;
  assign r = r_1; //(module output)
  /* fppow16.vhdl:2085:15  */
  assign cin_1_d1 = n1856; // (signal)
  /* fppow16.vhdl:2085:25  */
  assign cin_1_d2 = n1857; // (signal)
  /* fppow16.vhdl:2087:8  */
  assign x_1 = n1849; // (signal)
  /* fppow16.vhdl:2087:13  */
  assign x_1_d1 = n1858; // (signal)
  /* fppow16.vhdl:2089:8  */
  assign y_1 = n1851; // (signal)
  /* fppow16.vhdl:2089:13  */
  assign y_1_d1 = n1859; // (signal)
  /* fppow16.vhdl:2091:8  */
  assign s_1 = n1854; // (signal)
  /* fppow16.vhdl:2093:8  */
  assign r_1 = n1855; // (signal)
  /* fppow16.vhdl:2106:15  */
  assign n1849 = {1'b0, x};
  /* fppow16.vhdl:2107:15  */
  assign n1851 = {1'b0, y};
  /* fppow16.vhdl:2108:18  */
  assign n1852 = x_1_d1 + y_1_d1;
  /* fppow16.vhdl:2108:27  */
  assign n1853 = {21'b0, cin_1_d2};  //  uext
  /* fppow16.vhdl:2108:27  */
  assign n1854 = n1852 + n1853;
  /* fppow16.vhdl:2109:14  */
  assign n1855 = s_1[20:0]; // extract
  /* fppow16.vhdl:2098:10  */
  always @(posedge clk)
    n1856 <= cin_1;
  /* fppow16.vhdl:2098:10  */
  always @(posedge clk)
    n1857 <= cin_1_d1;
  /* fppow16.vhdl:2098:10  */
  always @(posedge clk)
    n1858 <= x_1;
  /* fppow16.vhdl:2098:10  */
  always @(posedge clk)
    n1859 <= y_1;
endmodule

module inva0table_freq500_uid15
  (input  [6:0] x,
   output [7:0] y);
  wire [7:0] y0;
  wire [7:0] y1;
  wire n1454;
  wire n1457;
  wire n1460;
  wire n1463;
  wire n1466;
  wire n1469;
  wire n1472;
  wire n1475;
  wire n1478;
  wire n1481;
  wire n1484;
  wire n1487;
  wire n1490;
  wire n1493;
  wire n1496;
  wire n1499;
  wire n1502;
  wire n1505;
  wire n1508;
  wire n1511;
  wire n1514;
  wire n1517;
  wire n1520;
  wire n1523;
  wire n1526;
  wire n1529;
  wire n1532;
  wire n1535;
  wire n1538;
  wire n1541;
  wire n1544;
  wire n1547;
  wire n1550;
  wire n1553;
  wire n1556;
  wire n1559;
  wire n1562;
  wire n1565;
  wire n1568;
  wire n1571;
  wire n1574;
  wire n1577;
  wire n1580;
  wire n1583;
  wire n1586;
  wire n1589;
  wire n1592;
  wire n1595;
  wire n1598;
  wire n1601;
  wire n1604;
  wire n1607;
  wire n1610;
  wire n1613;
  wire n1616;
  wire n1619;
  wire n1622;
  wire n1625;
  wire n1628;
  wire n1631;
  wire n1634;
  wire n1637;
  wire n1640;
  wire n1643;
  wire n1646;
  wire n1649;
  wire n1652;
  wire n1655;
  wire n1658;
  wire n1661;
  wire n1664;
  wire n1667;
  wire n1670;
  wire n1673;
  wire n1676;
  wire n1679;
  wire n1682;
  wire n1685;
  wire n1688;
  wire n1691;
  wire n1694;
  wire n1697;
  wire n1700;
  wire n1703;
  wire n1706;
  wire n1709;
  wire n1712;
  wire n1715;
  wire n1718;
  wire n1721;
  wire n1724;
  wire n1727;
  wire n1730;
  wire n1733;
  wire n1736;
  wire n1739;
  wire n1742;
  wire n1745;
  wire n1748;
  wire n1751;
  wire n1754;
  wire n1757;
  wire n1760;
  wire n1763;
  wire n1766;
  wire n1769;
  wire n1772;
  wire n1775;
  wire n1778;
  wire n1781;
  wire n1784;
  wire n1787;
  wire n1790;
  wire n1793;
  wire n1796;
  wire n1799;
  wire n1802;
  wire n1805;
  wire n1808;
  wire n1811;
  wire n1814;
  wire n1817;
  wire n1820;
  wire n1823;
  wire n1826;
  wire n1829;
  wire n1832;
  wire n1835;
  wire [127:0] n1837;
  reg [7:0] n1838;
  assign y = y1; //(module output)
  /* fppow16.vhdl:30:8  */
  assign y0 = n1838; // (signal)
  /* fppow16.vhdl:32:8  */
  assign y1 = y0; // (signal)
  /* fppow16.vhdl:36:18  */
  assign n1454 = x == 7'b0000000;
  /* fppow16.vhdl:37:18  */
  assign n1457 = x == 7'b0000001;
  /* fppow16.vhdl:38:18  */
  assign n1460 = x == 7'b0000010;
  /* fppow16.vhdl:39:18  */
  assign n1463 = x == 7'b0000011;
  /* fppow16.vhdl:40:18  */
  assign n1466 = x == 7'b0000100;
  /* fppow16.vhdl:41:18  */
  assign n1469 = x == 7'b0000101;
  /* fppow16.vhdl:42:18  */
  assign n1472 = x == 7'b0000110;
  /* fppow16.vhdl:43:18  */
  assign n1475 = x == 7'b0000111;
  /* fppow16.vhdl:44:18  */
  assign n1478 = x == 7'b0001000;
  /* fppow16.vhdl:45:18  */
  assign n1481 = x == 7'b0001001;
  /* fppow16.vhdl:46:18  */
  assign n1484 = x == 7'b0001010;
  /* fppow16.vhdl:47:18  */
  assign n1487 = x == 7'b0001011;
  /* fppow16.vhdl:48:18  */
  assign n1490 = x == 7'b0001100;
  /* fppow16.vhdl:49:18  */
  assign n1493 = x == 7'b0001101;
  /* fppow16.vhdl:50:18  */
  assign n1496 = x == 7'b0001110;
  /* fppow16.vhdl:51:18  */
  assign n1499 = x == 7'b0001111;
  /* fppow16.vhdl:52:18  */
  assign n1502 = x == 7'b0010000;
  /* fppow16.vhdl:53:18  */
  assign n1505 = x == 7'b0010001;
  /* fppow16.vhdl:54:18  */
  assign n1508 = x == 7'b0010010;
  /* fppow16.vhdl:55:18  */
  assign n1511 = x == 7'b0010011;
  /* fppow16.vhdl:56:18  */
  assign n1514 = x == 7'b0010100;
  /* fppow16.vhdl:57:18  */
  assign n1517 = x == 7'b0010101;
  /* fppow16.vhdl:58:18  */
  assign n1520 = x == 7'b0010110;
  /* fppow16.vhdl:59:18  */
  assign n1523 = x == 7'b0010111;
  /* fppow16.vhdl:60:18  */
  assign n1526 = x == 7'b0011000;
  /* fppow16.vhdl:61:18  */
  assign n1529 = x == 7'b0011001;
  /* fppow16.vhdl:62:18  */
  assign n1532 = x == 7'b0011010;
  /* fppow16.vhdl:63:18  */
  assign n1535 = x == 7'b0011011;
  /* fppow16.vhdl:64:18  */
  assign n1538 = x == 7'b0011100;
  /* fppow16.vhdl:65:18  */
  assign n1541 = x == 7'b0011101;
  /* fppow16.vhdl:66:18  */
  assign n1544 = x == 7'b0011110;
  /* fppow16.vhdl:67:18  */
  assign n1547 = x == 7'b0011111;
  /* fppow16.vhdl:68:18  */
  assign n1550 = x == 7'b0100000;
  /* fppow16.vhdl:69:18  */
  assign n1553 = x == 7'b0100001;
  /* fppow16.vhdl:70:18  */
  assign n1556 = x == 7'b0100010;
  /* fppow16.vhdl:71:18  */
  assign n1559 = x == 7'b0100011;
  /* fppow16.vhdl:72:18  */
  assign n1562 = x == 7'b0100100;
  /* fppow16.vhdl:73:18  */
  assign n1565 = x == 7'b0100101;
  /* fppow16.vhdl:74:18  */
  assign n1568 = x == 7'b0100110;
  /* fppow16.vhdl:75:18  */
  assign n1571 = x == 7'b0100111;
  /* fppow16.vhdl:76:18  */
  assign n1574 = x == 7'b0101000;
  /* fppow16.vhdl:77:18  */
  assign n1577 = x == 7'b0101001;
  /* fppow16.vhdl:78:18  */
  assign n1580 = x == 7'b0101010;
  /* fppow16.vhdl:79:18  */
  assign n1583 = x == 7'b0101011;
  /* fppow16.vhdl:80:18  */
  assign n1586 = x == 7'b0101100;
  /* fppow16.vhdl:81:18  */
  assign n1589 = x == 7'b0101101;
  /* fppow16.vhdl:82:18  */
  assign n1592 = x == 7'b0101110;
  /* fppow16.vhdl:83:18  */
  assign n1595 = x == 7'b0101111;
  /* fppow16.vhdl:84:18  */
  assign n1598 = x == 7'b0110000;
  /* fppow16.vhdl:85:18  */
  assign n1601 = x == 7'b0110001;
  /* fppow16.vhdl:86:18  */
  assign n1604 = x == 7'b0110010;
  /* fppow16.vhdl:87:18  */
  assign n1607 = x == 7'b0110011;
  /* fppow16.vhdl:88:18  */
  assign n1610 = x == 7'b0110100;
  /* fppow16.vhdl:89:18  */
  assign n1613 = x == 7'b0110101;
  /* fppow16.vhdl:90:18  */
  assign n1616 = x == 7'b0110110;
  /* fppow16.vhdl:91:18  */
  assign n1619 = x == 7'b0110111;
  /* fppow16.vhdl:92:18  */
  assign n1622 = x == 7'b0111000;
  /* fppow16.vhdl:93:18  */
  assign n1625 = x == 7'b0111001;
  /* fppow16.vhdl:94:18  */
  assign n1628 = x == 7'b0111010;
  /* fppow16.vhdl:95:18  */
  assign n1631 = x == 7'b0111011;
  /* fppow16.vhdl:96:18  */
  assign n1634 = x == 7'b0111100;
  /* fppow16.vhdl:97:18  */
  assign n1637 = x == 7'b0111101;
  /* fppow16.vhdl:98:18  */
  assign n1640 = x == 7'b0111110;
  /* fppow16.vhdl:99:18  */
  assign n1643 = x == 7'b0111111;
  /* fppow16.vhdl:100:18  */
  assign n1646 = x == 7'b1000000;
  /* fppow16.vhdl:101:18  */
  assign n1649 = x == 7'b1000001;
  /* fppow16.vhdl:102:18  */
  assign n1652 = x == 7'b1000010;
  /* fppow16.vhdl:103:18  */
  assign n1655 = x == 7'b1000011;
  /* fppow16.vhdl:104:18  */
  assign n1658 = x == 7'b1000100;
  /* fppow16.vhdl:105:18  */
  assign n1661 = x == 7'b1000101;
  /* fppow16.vhdl:106:18  */
  assign n1664 = x == 7'b1000110;
  /* fppow16.vhdl:107:18  */
  assign n1667 = x == 7'b1000111;
  /* fppow16.vhdl:108:18  */
  assign n1670 = x == 7'b1001000;
  /* fppow16.vhdl:109:18  */
  assign n1673 = x == 7'b1001001;
  /* fppow16.vhdl:110:18  */
  assign n1676 = x == 7'b1001010;
  /* fppow16.vhdl:111:18  */
  assign n1679 = x == 7'b1001011;
  /* fppow16.vhdl:112:18  */
  assign n1682 = x == 7'b1001100;
  /* fppow16.vhdl:113:18  */
  assign n1685 = x == 7'b1001101;
  /* fppow16.vhdl:114:18  */
  assign n1688 = x == 7'b1001110;
  /* fppow16.vhdl:115:18  */
  assign n1691 = x == 7'b1001111;
  /* fppow16.vhdl:116:18  */
  assign n1694 = x == 7'b1010000;
  /* fppow16.vhdl:117:18  */
  assign n1697 = x == 7'b1010001;
  /* fppow16.vhdl:118:18  */
  assign n1700 = x == 7'b1010010;
  /* fppow16.vhdl:119:18  */
  assign n1703 = x == 7'b1010011;
  /* fppow16.vhdl:120:18  */
  assign n1706 = x == 7'b1010100;
  /* fppow16.vhdl:121:18  */
  assign n1709 = x == 7'b1010101;
  /* fppow16.vhdl:122:18  */
  assign n1712 = x == 7'b1010110;
  /* fppow16.vhdl:123:18  */
  assign n1715 = x == 7'b1010111;
  /* fppow16.vhdl:124:18  */
  assign n1718 = x == 7'b1011000;
  /* fppow16.vhdl:125:18  */
  assign n1721 = x == 7'b1011001;
  /* fppow16.vhdl:126:18  */
  assign n1724 = x == 7'b1011010;
  /* fppow16.vhdl:127:18  */
  assign n1727 = x == 7'b1011011;
  /* fppow16.vhdl:128:18  */
  assign n1730 = x == 7'b1011100;
  /* fppow16.vhdl:129:18  */
  assign n1733 = x == 7'b1011101;
  /* fppow16.vhdl:130:18  */
  assign n1736 = x == 7'b1011110;
  /* fppow16.vhdl:131:18  */
  assign n1739 = x == 7'b1011111;
  /* fppow16.vhdl:132:18  */
  assign n1742 = x == 7'b1100000;
  /* fppow16.vhdl:133:18  */
  assign n1745 = x == 7'b1100001;
  /* fppow16.vhdl:134:18  */
  assign n1748 = x == 7'b1100010;
  /* fppow16.vhdl:135:18  */
  assign n1751 = x == 7'b1100011;
  /* fppow16.vhdl:136:18  */
  assign n1754 = x == 7'b1100100;
  /* fppow16.vhdl:137:18  */
  assign n1757 = x == 7'b1100101;
  /* fppow16.vhdl:138:18  */
  assign n1760 = x == 7'b1100110;
  /* fppow16.vhdl:139:18  */
  assign n1763 = x == 7'b1100111;
  /* fppow16.vhdl:140:18  */
  assign n1766 = x == 7'b1101000;
  /* fppow16.vhdl:141:18  */
  assign n1769 = x == 7'b1101001;
  /* fppow16.vhdl:142:18  */
  assign n1772 = x == 7'b1101010;
  /* fppow16.vhdl:143:18  */
  assign n1775 = x == 7'b1101011;
  /* fppow16.vhdl:144:18  */
  assign n1778 = x == 7'b1101100;
  /* fppow16.vhdl:145:18  */
  assign n1781 = x == 7'b1101101;
  /* fppow16.vhdl:146:18  */
  assign n1784 = x == 7'b1101110;
  /* fppow16.vhdl:147:18  */
  assign n1787 = x == 7'b1101111;
  /* fppow16.vhdl:148:18  */
  assign n1790 = x == 7'b1110000;
  /* fppow16.vhdl:149:18  */
  assign n1793 = x == 7'b1110001;
  /* fppow16.vhdl:150:18  */
  assign n1796 = x == 7'b1110010;
  /* fppow16.vhdl:151:18  */
  assign n1799 = x == 7'b1110011;
  /* fppow16.vhdl:152:18  */
  assign n1802 = x == 7'b1110100;
  /* fppow16.vhdl:153:18  */
  assign n1805 = x == 7'b1110101;
  /* fppow16.vhdl:154:18  */
  assign n1808 = x == 7'b1110110;
  /* fppow16.vhdl:155:18  */
  assign n1811 = x == 7'b1110111;
  /* fppow16.vhdl:156:18  */
  assign n1814 = x == 7'b1111000;
  /* fppow16.vhdl:157:18  */
  assign n1817 = x == 7'b1111001;
  /* fppow16.vhdl:158:18  */
  assign n1820 = x == 7'b1111010;
  /* fppow16.vhdl:159:18  */
  assign n1823 = x == 7'b1111011;
  /* fppow16.vhdl:160:18  */
  assign n1826 = x == 7'b1111100;
  /* fppow16.vhdl:161:18  */
  assign n1829 = x == 7'b1111101;
  /* fppow16.vhdl:162:18  */
  assign n1832 = x == 7'b1111110;
  /* fppow16.vhdl:163:18  */
  assign n1835 = x == 7'b1111111;
  assign n1837 = {n1835, n1832, n1829, n1826, n1823, n1820, n1817, n1814, n1811, n1808, n1805, n1802, n1799, n1796, n1793, n1790, n1787, n1784, n1781, n1778, n1775, n1772, n1769, n1766, n1763, n1760, n1757, n1754, n1751, n1748, n1745, n1742, n1739, n1736, n1733, n1730, n1727, n1724, n1721, n1718, n1715, n1712, n1709, n1706, n1703, n1700, n1697, n1694, n1691, n1688, n1685, n1682, n1679, n1676, n1673, n1670, n1667, n1664, n1661, n1658, n1655, n1652, n1649, n1646, n1643, n1640, n1637, n1634, n1631, n1628, n1625, n1622, n1619, n1616, n1613, n1610, n1607, n1604, n1601, n1598, n1595, n1592, n1589, n1586, n1583, n1580, n1577, n1574, n1571, n1568, n1565, n1562, n1559, n1556, n1553, n1550, n1547, n1544, n1541, n1538, n1535, n1532, n1529, n1526, n1523, n1520, n1517, n1514, n1511, n1508, n1505, n1502, n1499, n1496, n1493, n1490, n1487, n1484, n1481, n1478, n1475, n1472, n1469, n1466, n1463, n1460, n1457, n1454};
  /* fppow16.vhdl:35:4  */
  always @*
    case (n1837)
      128'b10000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1838 = 8'b10000001;
      128'b01000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1838 = 8'b10000010;
      128'b00100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1838 = 8'b10000010;
      128'b00010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1838 = 8'b10000011;
      128'b00001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1838 = 8'b10000011;
      128'b00000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1838 = 8'b10000100;
      128'b00000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1838 = 8'b10000100;
      128'b00000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1838 = 8'b10000101;
      128'b00000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1838 = 8'b10000101;
      128'b00000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1838 = 8'b10000110;
      128'b00000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1838 = 8'b10000110;
      128'b00000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1838 = 8'b10000111;
      128'b00000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1838 = 8'b10000111;
      128'b00000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1838 = 8'b10001000;
      128'b00000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1838 = 8'b10001000;
      128'b00000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1838 = 8'b10001001;
      128'b00000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1838 = 8'b10001010;
      128'b00000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1838 = 8'b10001010;
      128'b00000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1838 = 8'b10001011;
      128'b00000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1838 = 8'b10001011;
      128'b00000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1838 = 8'b10001100;
      128'b00000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1838 = 8'b10001101;
      128'b00000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1838 = 8'b10001101;
      128'b00000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1838 = 8'b10001110;
      128'b00000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1838 = 8'b10001110;
      128'b00000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1838 = 8'b10001111;
      128'b00000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1838 = 8'b10010000;
      128'b00000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1838 = 8'b10010000;
      128'b00000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1838 = 8'b10010001;
      128'b00000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1838 = 8'b10010001;
      128'b00000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1838 = 8'b10010010;
      128'b00000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1838 = 8'b10010011;
      128'b00000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1838 = 8'b10010011;
      128'b00000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1838 = 8'b10010100;
      128'b00000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1838 = 8'b10010101;
      128'b00000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1838 = 8'b10010101;
      128'b00000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1838 = 8'b10010110;
      128'b00000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1838 = 8'b10010111;
      128'b00000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1838 = 8'b10011000;
      128'b00000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1838 = 8'b10011000;
      128'b00000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1838 = 8'b10011001;
      128'b00000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1838 = 8'b10011010;
      128'b00000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1838 = 8'b10011010;
      128'b00000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1838 = 8'b10011011;
      128'b00000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1838 = 8'b10011100;
      128'b00000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1838 = 8'b10011101;
      128'b00000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1838 = 8'b10011101;
      128'b00000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000: n1838 = 8'b10011110;
      128'b00000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000: n1838 = 8'b10011111;
      128'b00000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000: n1838 = 8'b10100000;
      128'b00000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000: n1838 = 8'b10100000;
      128'b00000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000: n1838 = 8'b10100001;
      128'b00000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000: n1838 = 8'b10100010;
      128'b00000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000: n1838 = 8'b10100011;
      128'b00000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000: n1838 = 8'b10100100;
      128'b00000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000: n1838 = 8'b10100100;
      128'b00000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000: n1838 = 8'b10100101;
      128'b00000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000: n1838 = 8'b10100110;
      128'b00000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000: n1838 = 8'b10100111;
      128'b00000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000: n1838 = 8'b10101000;
      128'b00000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000: n1838 = 8'b10101001;
      128'b00000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000: n1838 = 8'b10101001;
      128'b00000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000: n1838 = 8'b10101010;
      128'b00000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000: n1838 = 8'b10101011;
      128'b00000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000: n1838 = 8'b01010110;
      128'b00000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000: n1838 = 8'b01010111;
      128'b00000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000: n1838 = 8'b01010111;
      128'b00000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000: n1838 = 8'b01011000;
      128'b00000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000: n1838 = 8'b01011000;
      128'b00000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000: n1838 = 8'b01011001;
      128'b00000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000: n1838 = 8'b01011001;
      128'b00000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000: n1838 = 8'b01011010;
      128'b00000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000: n1838 = 8'b01011010;
      128'b00000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000: n1838 = 8'b01011011;
      128'b00000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000: n1838 = 8'b01011011;
      128'b00000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000: n1838 = 8'b01011100;
      128'b00000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000: n1838 = 8'b01011100;
      128'b00000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000: n1838 = 8'b01011101;
      128'b00000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000: n1838 = 8'b01011101;
      128'b00000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000: n1838 = 8'b01011110;
      128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000: n1838 = 8'b01011110;
      128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000: n1838 = 8'b01011111;
      128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000: n1838 = 8'b01011111;
      128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000: n1838 = 8'b01100000;
      128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000: n1838 = 8'b01100000;
      128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000: n1838 = 8'b01100001;
      128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000: n1838 = 8'b01100001;
      128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000: n1838 = 8'b01100010;
      128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000: n1838 = 8'b01100011;
      128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000: n1838 = 8'b01100011;
      128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000: n1838 = 8'b01100100;
      128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000: n1838 = 8'b01100100;
      128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000: n1838 = 8'b01100101;
      128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000: n1838 = 8'b01100110;
      128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000: n1838 = 8'b01100110;
      128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000: n1838 = 8'b01100111;
      128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000: n1838 = 8'b01101000;
      128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000: n1838 = 8'b01101000;
      128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000: n1838 = 8'b01101001;
      128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000: n1838 = 8'b01101010;
      128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000: n1838 = 8'b01101010;
      128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000: n1838 = 8'b01101011;
      128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000: n1838 = 8'b01101100;
      128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000: n1838 = 8'b01101100;
      128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000: n1838 = 8'b01101101;
      128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000: n1838 = 8'b01101110;
      128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000: n1838 = 8'b01101110;
      128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000: n1838 = 8'b01101111;
      128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000: n1838 = 8'b01110000;
      128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000: n1838 = 8'b01110001;
      128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000: n1838 = 8'b01110001;
      128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000: n1838 = 8'b01110010;
      128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000: n1838 = 8'b01110011;
      128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000: n1838 = 8'b01110100;
      128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000: n1838 = 8'b01110101;
      128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000: n1838 = 8'b01110110;
      128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000: n1838 = 8'b01110110;
      128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000: n1838 = 8'b01110111;
      128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000: n1838 = 8'b01111000;
      128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000: n1838 = 8'b01111001;
      128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000: n1838 = 8'b01111010;
      128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000: n1838 = 8'b01111011;
      128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000: n1838 = 8'b01111100;
      128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000: n1838 = 8'b01111101;
      128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000: n1838 = 8'b01111110;
      128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100: n1838 = 8'b01111111;
      128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010: n1838 = 8'b10000000;
      128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001: n1838 = 8'b10000000;
      default: n1838 = 8'bX;
    endcase
endmodule

module leftshifter10_by_max_10_freq500_uid13
  (input  clk,
   input  [9:0] x,
   input  [3:0] s,
   output [19:0] r);
  wire [3:0] ps;
  wire [3:0] ps_d1;
  wire [9:0] level0;
  wire [9:0] level0_d1;
  wire [9:0] level0_d2;
  wire [9:0] level0_d3;
  wire [10:0] level1;
  wire [10:0] level1_d1;
  wire [12:0] level2;
  wire [16:0] level3;
  wire [24:0] level4;
  wire [10:0] n1422;
  wire n1423;
  wire [10:0] n1424;
  wire [10:0] n1426;
  wire [12:0] n1428;
  wire n1429;
  wire [12:0] n1430;
  wire [12:0] n1432;
  wire [16:0] n1434;
  wire n1435;
  wire [16:0] n1436;
  wire [16:0] n1438;
  wire [24:0] n1440;
  wire n1441;
  wire [24:0] n1442;
  wire [24:0] n1444;
  wire [19:0] n1445;
  reg [3:0] n1446;
  reg [9:0] n1447;
  reg [9:0] n1448;
  reg [9:0] n1449;
  reg [10:0] n1450;
  assign r = n1445; //(module output)
  /* fppow16.vhdl:2021:12  */
  assign ps_d1 = n1446; // (signal)
  /* fppow16.vhdl:2023:16  */
  assign level0_d1 = n1447; // (signal)
  /* fppow16.vhdl:2023:27  */
  assign level0_d2 = n1448; // (signal)
  /* fppow16.vhdl:2023:38  */
  assign level0_d3 = n1449; // (signal)
  /* fppow16.vhdl:2025:8  */
  assign level1 = n1424; // (signal)
  /* fppow16.vhdl:2025:16  */
  assign level1_d1 = n1450; // (signal)
  /* fppow16.vhdl:2027:8  */
  assign level2 = n1430; // (signal)
  /* fppow16.vhdl:2029:8  */
  assign level3 = n1436; // (signal)
  /* fppow16.vhdl:2031:8  */
  assign level4 = n1442; // (signal)
  /* fppow16.vhdl:2046:23  */
  assign n1422 = {level0_d3, 1'b0};
  /* fppow16.vhdl:2046:52  */
  assign n1423 = ps[0]; // extract
  /* fppow16.vhdl:2046:45  */
  assign n1424 = n1423 ? n1422 : n1426;
  /* fppow16.vhdl:2046:90  */
  assign n1426 = {1'b0, level0_d3};
  /* fppow16.vhdl:2047:23  */
  assign n1428 = {level1_d1, 2'b00};
  /* fppow16.vhdl:2047:55  */
  assign n1429 = ps_d1[1]; // extract
  /* fppow16.vhdl:2047:45  */
  assign n1430 = n1429 ? n1428 : n1432;
  /* fppow16.vhdl:2047:93  */
  assign n1432 = {2'b00, level1_d1};
  /* fppow16.vhdl:2048:20  */
  assign n1434 = {level2, 4'b0000};
  /* fppow16.vhdl:2048:52  */
  assign n1435 = ps_d1[2]; // extract
  /* fppow16.vhdl:2048:42  */
  assign n1436 = n1435 ? n1434 : n1438;
  /* fppow16.vhdl:2048:90  */
  assign n1438 = {4'b0000, level2};
  /* fppow16.vhdl:2049:20  */
  assign n1440 = {level3, 8'b00000000};
  /* fppow16.vhdl:2049:52  */
  assign n1441 = ps_d1[3]; // extract
  /* fppow16.vhdl:2049:42  */
  assign n1442 = n1441 ? n1440 : n1444;
  /* fppow16.vhdl:2049:90  */
  assign n1444 = {8'b00000000, level3};
  /* fppow16.vhdl:2050:15  */
  assign n1445 = level4[19:0]; // extract
  /* fppow16.vhdl:2036:10  */
  always @(posedge clk)
    n1446 <= ps;
  /* fppow16.vhdl:2036:10  */
  always @(posedge clk)
    n1447 <= level0;
  /* fppow16.vhdl:2036:10  */
  always @(posedge clk)
    n1448 <= level0_d1;
  /* fppow16.vhdl:2036:10  */
  always @(posedge clk)
    n1449 <= level0_d2;
  /* fppow16.vhdl:2036:10  */
  always @(posedge clk)
    n1450 <= level1;
endmodule

module lzoc_17_freq500_uid11
  (input  clk,
   input  [16:0] i,
   input  ozb,
   output [4:0] o);
  wire sozb;
  wire sozb_d1;
  wire sozb_d2;
  wire [30:0] level5;
  wire [30:0] level5_d1;
  wire digit4;
  wire digit4_d1;
  wire digit4_d2;
  wire [14:0] level4;
  wire [14:0] level4_d1;
  wire digit3;
  wire digit3_d1;
  wire [6:0] level3;
  wire digit2;
  wire [2:0] level2;
  wire [2:0] level2_d1;
  wire [2:0] z;
  wire [1:0] lowbits;
  wire [2:0] outhighbits;
  wire [2:0] outhighbits_d1;
  wire ozb_d1;
  wire ozb_d2;
  wire ozb_d3;
  wire n1324;
  wire n1325;
  wire n1326;
  wire n1327;
  wire n1328;
  wire n1329;
  wire n1330;
  wire n1331;
  wire n1332;
  wire n1333;
  wire n1334;
  wire n1335;
  wire n1336;
  wire n1337;
  wire [3:0] n1338;
  wire [3:0] n1339;
  wire [3:0] n1340;
  wire [1:0] n1341;
  wire [13:0] n1342;
  wire [30:0] n1343;
  wire [15:0] n1345;
  wire [3:0] n1346;
  wire [3:0] n1347;
  wire [3:0] n1348;
  wire [3:0] n1349;
  wire [15:0] n1350;
  wire n1351;
  wire n1352;
  wire [14:0] n1354;
  wire [14:0] n1355;
  wire [14:0] n1356;
  wire [7:0] n1358;
  wire [3:0] n1359;
  wire [3:0] n1360;
  wire [7:0] n1361;
  wire n1362;
  wire n1363;
  wire [6:0] n1365;
  wire [6:0] n1366;
  wire [6:0] n1367;
  wire [3:0] n1369;
  wire [3:0] n1370;
  wire n1371;
  wire n1372;
  wire [2:0] n1374;
  wire [2:0] n1375;
  wire [2:0] n1376;
  wire n1377;
  wire [2:0] n1378;
  wire [2:0] n1379;
  wire n1382;
  wire n1385;
  wire n1388;
  wire n1391;
  wire [3:0] n1393;
  reg [1:0] n1394;
  wire [1:0] n1395;
  wire [2:0] n1396;
  wire [4:0] n1398;
  reg n1399;
  reg n1400;
  reg [30:0] n1401;
  reg n1402;
  reg n1403;
  reg [14:0] n1404;
  reg n1405;
  reg [2:0] n1406;
  reg [2:0] n1407;
  reg n1408;
  reg n1409;
  reg n1410;
  assign o = n1398; //(module output)
  /* fppow16.vhdl:1926:8  */
  assign sozb = ozb; // (signal)
  /* fppow16.vhdl:1926:14  */
  assign sozb_d1 = n1399; // (signal)
  /* fppow16.vhdl:1926:23  */
  assign sozb_d2 = n1400; // (signal)
  /* fppow16.vhdl:1928:8  */
  assign level5 = n1343; // (signal)
  /* fppow16.vhdl:1928:16  */
  assign level5_d1 = n1401; // (signal)
  /* fppow16.vhdl:1930:8  */
  assign digit4 = n1352; // (signal)
  /* fppow16.vhdl:1930:16  */
  assign digit4_d1 = n1402; // (signal)
  /* fppow16.vhdl:1930:27  */
  assign digit4_d2 = n1403; // (signal)
  /* fppow16.vhdl:1932:8  */
  assign level4 = n1355; // (signal)
  /* fppow16.vhdl:1932:16  */
  assign level4_d1 = n1404; // (signal)
  /* fppow16.vhdl:1934:8  */
  assign digit3 = n1363; // (signal)
  /* fppow16.vhdl:1934:16  */
  assign digit3_d1 = n1405; // (signal)
  /* fppow16.vhdl:1936:8  */
  assign level3 = n1366; // (signal)
  /* fppow16.vhdl:1938:8  */
  assign digit2 = n1372; // (signal)
  /* fppow16.vhdl:1940:8  */
  assign level2 = n1375; // (signal)
  /* fppow16.vhdl:1940:16  */
  assign level2_d1 = n1406; // (signal)
  /* fppow16.vhdl:1942:8  */
  assign z = n1378; // (signal)
  /* fppow16.vhdl:1944:8  */
  assign lowbits = n1394; // (signal)
  /* fppow16.vhdl:1946:8  */
  assign outhighbits = n1396; // (signal)
  /* fppow16.vhdl:1946:21  */
  assign outhighbits_d1 = n1407; // (signal)
  /* fppow16.vhdl:1948:8  */
  assign ozb_d1 = n1408; // (signal)
  /* fppow16.vhdl:1948:16  */
  assign ozb_d2 = n1409; // (signal)
  /* fppow16.vhdl:1948:24  */
  assign ozb_d3 = n1410; // (signal)
  /* fppow16.vhdl:1970:34  */
  assign n1324 = ~sozb;
  /* fppow16.vhdl:1970:34  */
  assign n1325 = ~sozb;
  /* fppow16.vhdl:1970:34  */
  assign n1326 = ~sozb;
  /* fppow16.vhdl:1970:34  */
  assign n1327 = ~sozb;
  /* fppow16.vhdl:1970:34  */
  assign n1328 = ~sozb;
  /* fppow16.vhdl:1970:34  */
  assign n1329 = ~sozb;
  /* fppow16.vhdl:1970:34  */
  assign n1330 = ~sozb;
  /* fppow16.vhdl:1970:34  */
  assign n1331 = ~sozb;
  /* fppow16.vhdl:1970:34  */
  assign n1332 = ~sozb;
  /* fppow16.vhdl:1970:34  */
  assign n1333 = ~sozb;
  /* fppow16.vhdl:1970:34  */
  assign n1334 = ~sozb;
  /* fppow16.vhdl:1970:34  */
  assign n1335 = ~sozb;
  /* fppow16.vhdl:1970:34  */
  assign n1336 = ~sozb;
  /* fppow16.vhdl:1970:34  */
  assign n1337 = ~sozb;
  assign n1338 = {n1337, n1336, n1335, n1334};
  assign n1339 = {n1333, n1332, n1331, n1330};
  assign n1340 = {n1329, n1328, n1327, n1326};
  assign n1341 = {n1325, n1324};
  assign n1342 = {n1338, n1339, n1340, n1341};
  /* fppow16.vhdl:1970:16  */
  assign n1343 = {i, n1342};
  /* fppow16.vhdl:1972:28  */
  assign n1345 = level5[30:15]; // extract
  assign n1346 = {sozb, sozb, sozb, sozb};
  assign n1347 = {sozb, sozb, sozb, sozb};
  assign n1348 = {sozb, sozb, sozb, sozb};
  assign n1349 = {sozb, sozb, sozb, sozb};
  assign n1350 = {n1346, n1347, n1348, n1349};
  /* fppow16.vhdl:1972:43  */
  assign n1351 = n1345 == n1350;
  /* fppow16.vhdl:1972:17  */
  assign n1352 = n1351 ? 1'b1 : 1'b0;
  /* fppow16.vhdl:1973:22  */
  assign n1354 = level5_d1[14:0]; // extract
  /* fppow16.vhdl:1973:36  */
  assign n1355 = digit4_d1 ? n1354 : n1356;
  /* fppow16.vhdl:1973:69  */
  assign n1356 = level5_d1[30:16]; // extract
  /* fppow16.vhdl:1974:28  */
  assign n1358 = level4[14:7]; // extract
  assign n1359 = {sozb_d1, sozb_d1, sozb_d1, sozb_d1};
  assign n1360 = {sozb_d1, sozb_d1, sozb_d1, sozb_d1};
  assign n1361 = {n1359, n1360};
  /* fppow16.vhdl:1974:42  */
  assign n1362 = n1358 == n1361;
  /* fppow16.vhdl:1974:17  */
  assign n1363 = n1362 ? 1'b1 : 1'b0;
  /* fppow16.vhdl:1975:22  */
  assign n1365 = level4_d1[6:0]; // extract
  /* fppow16.vhdl:1975:35  */
  assign n1366 = digit3_d1 ? n1365 : n1367;
  /* fppow16.vhdl:1975:68  */
  assign n1367 = level4_d1[14:8]; // extract
  /* fppow16.vhdl:1976:28  */
  assign n1369 = level3[6:3]; // extract
  assign n1370 = {sozb_d2, sozb_d2, sozb_d2, sozb_d2};
  /* fppow16.vhdl:1976:41  */
  assign n1371 = n1369 == n1370;
  /* fppow16.vhdl:1976:17  */
  assign n1372 = n1371 ? 1'b1 : 1'b0;
  /* fppow16.vhdl:1977:19  */
  assign n1374 = level3[2:0]; // extract
  /* fppow16.vhdl:1977:32  */
  assign n1375 = digit2 ? n1374 : n1376;
  /* fppow16.vhdl:1977:59  */
  assign n1376 = level3[6:4]; // extract
  /* fppow16.vhdl:1979:30  */
  assign n1377 = ~ozb_d3;
  /* fppow16.vhdl:1979:19  */
  assign n1378 = n1377 ? level2_d1 : n1379;
  /* fppow16.vhdl:1979:41  */
  assign n1379 = ~level2_d1;
  /* fppow16.vhdl:1981:12  */
  assign n1382 = z == 3'b000;
  /* fppow16.vhdl:1982:12  */
  assign n1385 = z == 3'b001;
  /* fppow16.vhdl:1983:12  */
  assign n1388 = z == 3'b010;
  /* fppow16.vhdl:1984:12  */
  assign n1391 = z == 3'b011;
  assign n1393 = {n1391, n1388, n1385, n1382};
  /* fppow16.vhdl:1980:4  */
  always @*
    case (n1393)
      4'b1000: n1394 = 2'b01;
      4'b0100: n1394 = 2'b01;
      4'b0010: n1394 = 2'b10;
      4'b0001: n1394 = 2'b11;
      default: n1394 = 2'b00;
    endcase
  /* fppow16.vhdl:1986:29  */
  assign n1395 = {digit4_d2, digit3_d1};
  /* fppow16.vhdl:1986:50  */
  assign n1396 = {n1395, digit2};
  /* fppow16.vhdl:1987:24  */
  assign n1398 = {outhighbits_d1, lowbits};
  /* fppow16.vhdl:1953:10  */
  always @(posedge clk)
    n1399 <= sozb;
  /* fppow16.vhdl:1953:10  */
  always @(posedge clk)
    n1400 <= sozb_d1;
  /* fppow16.vhdl:1953:10  */
  always @(posedge clk)
    n1401 <= level5;
  /* fppow16.vhdl:1953:10  */
  always @(posedge clk)
    n1402 <= digit4;
  /* fppow16.vhdl:1953:10  */
  always @(posedge clk)
    n1403 <= digit4_d1;
  /* fppow16.vhdl:1953:10  */
  always @(posedge clk)
    n1404 <= level4;
  /* fppow16.vhdl:1953:10  */
  always @(posedge clk)
    n1405 <= digit3;
  /* fppow16.vhdl:1953:10  */
  always @(posedge clk)
    n1406 <= level2;
  /* fppow16.vhdl:1953:10  */
  always @(posedge clk)
    n1407 <= outhighbits;
  /* fppow16.vhdl:1953:10  */
  always @(posedge clk)
    n1408 <= ozb;
  /* fppow16.vhdl:1953:10  */
  always @(posedge clk)
    n1409 <= ozb_d1;
  /* fppow16.vhdl:1953:10  */
  always @(posedge clk)
    n1410 <= ozb_d2;
endmodule

module fpexp_5_10_freq500_uid66
  (input  clk,
   input  [25:0] x,
   output [17:0] r);
  wire [1:0] xexn;
  wire [1:0] xexn_d1;
  wire [1:0] xexn_d2;
  wire [1:0] xexn_d3;
  wire [1:0] xexn_d4;
  wire [1:0] xexn_d5;
  wire [1:0] xexn_d6;
  wire xsign;
  wire xsign_d1;
  wire xsign_d2;
  wire xsign_d3;
  wire xsign_d4;
  wire xsign_d5;
  wire xsign_d6;
  wire [4:0] xexpfield;
  wire [4:0] xexpfield_d1;
  wire [17:0] xfrac;
  wire [6:0] e0;
  wire [6:0] e0_d1;
  wire [6:0] e0_d2;
  wire [6:0] e0_d3;
  wire [6:0] e0_d4;
  wire [6:0] e0_d5;
  wire [6:0] e0_d6;
  wire [6:0] e0_d7;
  wire [6:0] e0_d8;
  wire [6:0] e0_d9;
  wire [6:0] e0_d10;
  wire [6:0] e0_d11;
  wire [6:0] e0_d12;
  wire [6:0] e0_d13;
  wire [6:0] shiftval;
  wire resultwillbeone;
  wire resultwillbeone_d1;
  wire [18:0] mxu;
  wire [5:0] maxshift;
  wire [5:0] maxshift_d1;
  wire [5:0] maxshift_d2;
  wire [5:0] maxshift_d3;
  wire [5:0] maxshift_d4;
  wire [5:0] maxshift_d5;
  wire [5:0] maxshift_d6;
  wire [5:0] maxshift_d7;
  wire [5:0] maxshift_d8;
  wire [5:0] maxshift_d9;
  wire [5:0] maxshift_d10;
  wire [5:0] maxshift_d11;
  wire [5:0] maxshift_d12;
  wire [5:0] maxshift_d13;
  wire overflow0;
  wire [4:0] shiftvalin;
  wire [34:0] fixx0;
  wire [16:0] ufixx;
  wire [13:0] expy;
  wire [5:0] k;
  wire [5:0] k_d1;
  wire [5:0] k_d2;
  wire neednonorm;
  wire [16:0] preroundbiassig;
  wire roundbit;
  wire [16:0] roundnormaddend;
  wire [16:0] roundedexpsigres;
  wire [16:0] roundedexpsig;
  wire ofl1;
  wire ofl1_d1;
  wire ofl1_d2;
  wire ofl1_d3;
  wire ofl1_d4;
  wire ofl1_d5;
  wire ofl2;
  wire ofl3;
  wire ofl3_d1;
  wire ofl3_d2;
  wire ofl3_d3;
  wire ofl3_d4;
  wire ofl3_d5;
  wire ofl3_d6;
  wire ofl;
  wire ufl1;
  wire ufl2;
  wire ufl2_d1;
  wire ufl2_d2;
  wire ufl2_d3;
  wire ufl2_d4;
  wire ufl2_d5;
  wire ufl2_d6;
  wire ufl3;
  wire ufl3_d1;
  wire ufl3_d2;
  wire ufl3_d3;
  wire ufl3_d4;
  wire ufl3_d5;
  wire ufl;
  wire [1:0] rexn;
  wire [1:0] n1127;
  wire n1128;
  wire [4:0] n1129;
  wire [17:0] n1130;
  wire [6:0] n1133;
  wire [6:0] n1134;
  wire n1135;
  wire [18:0] n1137;
  wire n1139;
  wire n1140;
  wire [5:0] n1141;
  wire n1142;
  wire n1143;
  wire [4:0] n1145;
  wire [34:0] mantissa_shift_n1146;
  wire [16:0] n1149;
  wire n1150;
  wire [16:0] n1151;
  wire [13:0] exp_helper_n1153;
  wire [5:0] exp_helper_n1154;
  wire n1159;
  wire [9:0] n1160;
  wire [16:0] n1162;
  wire [16:0] n1163;
  wire [9:0] n1164;
  wire [16:0] n1166;
  wire n1167;
  wire n1168;
  wire n1169;
  wire n1170;
  wire [6:0] n1171;
  wire [15:0] n1173;
  wire [16:0] n1174;
  localparam n1175 = 1'b0;
  wire [16:0] roundedexpsigoperandadder_n1176;
  wire n1180;
  wire [16:0] n1181;
  wire n1183;
  wire n1184;
  wire n1185;
  wire n1186;
  wire n1187;
  wire n1188;
  wire n1189;
  wire n1190;
  wire n1191;
  wire n1192;
  wire n1193;
  wire n1194;
  wire n1195;
  wire n1196;
  wire n1197;
  wire n1198;
  wire n1199;
  wire n1200;
  wire n1201;
  wire n1202;
  wire n1203;
  wire n1204;
  wire n1205;
  wire n1206;
  wire n1207;
  wire n1208;
  wire n1209;
  wire n1210;
  wire n1211;
  wire n1212;
  wire n1213;
  wire n1214;
  wire n1215;
  wire n1216;
  wire n1217;
  wire n1218;
  wire n1219;
  wire n1220;
  wire n1221;
  wire n1222;
  wire n1223;
  wire n1224;
  wire n1225;
  wire n1226;
  wire n1227;
  wire n1228;
  wire n1229;
  wire n1232;
  wire [1:0] n1233;
  wire [1:0] n1235;
  wire [1:0] n1237;
  wire [2:0] n1240;
  wire [14:0] n1241;
  wire [17:0] n1242;
  reg [1:0] n1243;
  reg [1:0] n1244;
  reg [1:0] n1245;
  reg [1:0] n1246;
  reg [1:0] n1247;
  reg [1:0] n1248;
  reg n1249;
  reg n1250;
  reg n1251;
  reg n1252;
  reg n1253;
  reg n1254;
  reg [4:0] n1255;
  reg [6:0] n1256;
  reg [6:0] n1257;
  reg [6:0] n1258;
  reg [6:0] n1259;
  reg [6:0] n1260;
  reg [6:0] n1261;
  reg [6:0] n1262;
  reg [6:0] n1263;
  reg [6:0] n1264;
  reg [6:0] n1265;
  reg [6:0] n1266;
  reg [6:0] n1267;
  reg [6:0] n1268;
  reg n1269;
  reg [5:0] n1270;
  reg [5:0] n1271;
  reg [5:0] n1272;
  reg [5:0] n1273;
  reg [5:0] n1274;
  reg [5:0] n1275;
  reg [5:0] n1276;
  reg [5:0] n1277;
  reg [5:0] n1278;
  reg [5:0] n1279;
  reg [5:0] n1280;
  reg [5:0] n1281;
  reg [5:0] n1282;
  reg [5:0] n1283;
  reg [5:0] n1284;
  reg n1285;
  reg n1286;
  reg n1287;
  reg n1288;
  reg n1289;
  reg n1290;
  reg n1291;
  reg n1292;
  reg n1293;
  reg n1294;
  reg n1295;
  reg n1296;
  reg n1297;
  reg n1298;
  reg n1299;
  reg n1300;
  reg n1301;
  reg n1302;
  reg n1303;
  reg n1304;
  reg n1305;
  reg n1306;
  assign r = n1242; //(module output)
  /* fppow16.vhdl:4667:8  */
  assign xexn = n1127; // (signal)
  /* fppow16.vhdl:4667:14  */
  assign xexn_d1 = n1243; // (signal)
  /* fppow16.vhdl:4667:23  */
  assign xexn_d2 = n1244; // (signal)
  /* fppow16.vhdl:4667:32  */
  assign xexn_d3 = n1245; // (signal)
  /* fppow16.vhdl:4667:41  */
  assign xexn_d4 = n1246; // (signal)
  /* fppow16.vhdl:4667:50  */
  assign xexn_d5 = n1247; // (signal)
  /* fppow16.vhdl:4667:59  */
  assign xexn_d6 = n1248; // (signal)
  /* fppow16.vhdl:4669:8  */
  assign xsign = n1128; // (signal)
  /* fppow16.vhdl:4669:15  */
  assign xsign_d1 = n1249; // (signal)
  /* fppow16.vhdl:4669:25  */
  assign xsign_d2 = n1250; // (signal)
  /* fppow16.vhdl:4669:35  */
  assign xsign_d3 = n1251; // (signal)
  /* fppow16.vhdl:4669:45  */
  assign xsign_d4 = n1252; // (signal)
  /* fppow16.vhdl:4669:55  */
  assign xsign_d5 = n1253; // (signal)
  /* fppow16.vhdl:4669:65  */
  assign xsign_d6 = n1254; // (signal)
  /* fppow16.vhdl:4671:8  */
  assign xexpfield = n1129; // (signal)
  /* fppow16.vhdl:4671:19  */
  assign xexpfield_d1 = n1255; // (signal)
  /* fppow16.vhdl:4673:8  */
  assign xfrac = n1130; // (signal)
  /* fppow16.vhdl:4675:8  */
  assign e0 = 7'b0000010; // (signal)
  /* fppow16.vhdl:4675:12  */
  assign e0_d1 = n1256; // (signal)
  /* fppow16.vhdl:4675:19  */
  assign e0_d2 = n1257; // (signal)
  /* fppow16.vhdl:4675:26  */
  assign e0_d3 = n1258; // (signal)
  /* fppow16.vhdl:4675:33  */
  assign e0_d4 = n1259; // (signal)
  /* fppow16.vhdl:4675:40  */
  assign e0_d5 = n1260; // (signal)
  /* fppow16.vhdl:4675:47  */
  assign e0_d6 = n1261; // (signal)
  /* fppow16.vhdl:4675:54  */
  assign e0_d7 = n1262; // (signal)
  /* fppow16.vhdl:4675:61  */
  assign e0_d8 = n1263; // (signal)
  /* fppow16.vhdl:4675:68  */
  assign e0_d9 = n1264; // (signal)
  /* fppow16.vhdl:4675:75  */
  assign e0_d10 = n1265; // (signal)
  /* fppow16.vhdl:4675:83  */
  assign e0_d11 = n1266; // (signal)
  /* fppow16.vhdl:4675:91  */
  assign e0_d12 = n1267; // (signal)
  /* fppow16.vhdl:4675:99  */
  assign e0_d13 = n1268; // (signal)
  /* fppow16.vhdl:4677:8  */
  assign shiftval = n1134; // (signal)
  /* fppow16.vhdl:4679:8  */
  assign resultwillbeone = n1135; // (signal)
  /* fppow16.vhdl:4679:25  */
  assign resultwillbeone_d1 = n1269; // (signal)
  /* fppow16.vhdl:4681:8  */
  assign mxu = n1137; // (signal)
  /* fppow16.vhdl:4683:8  */
  assign maxshift = 6'b010000; // (signal)
  /* fppow16.vhdl:4683:18  */
  assign maxshift_d1 = n1270; // (signal)
  /* fppow16.vhdl:4683:31  */
  assign maxshift_d2 = n1271; // (signal)
  /* fppow16.vhdl:4683:44  */
  assign maxshift_d3 = n1272; // (signal)
  /* fppow16.vhdl:4683:57  */
  assign maxshift_d4 = n1273; // (signal)
  /* fppow16.vhdl:4683:70  */
  assign maxshift_d5 = n1274; // (signal)
  /* fppow16.vhdl:4683:83  */
  assign maxshift_d6 = n1275; // (signal)
  /* fppow16.vhdl:4683:96  */
  assign maxshift_d7 = n1276; // (signal)
  /* fppow16.vhdl:4683:109  */
  assign maxshift_d8 = n1277; // (signal)
  /* fppow16.vhdl:4683:122  */
  assign maxshift_d9 = n1278; // (signal)
  /* fppow16.vhdl:4683:135  */
  assign maxshift_d10 = n1279; // (signal)
  /* fppow16.vhdl:4683:149  */
  assign maxshift_d11 = n1280; // (signal)
  /* fppow16.vhdl:4683:163  */
  assign maxshift_d12 = n1281; // (signal)
  /* fppow16.vhdl:4683:177  */
  assign maxshift_d13 = n1282; // (signal)
  /* fppow16.vhdl:4685:8  */
  assign overflow0 = n1143; // (signal)
  /* fppow16.vhdl:4687:8  */
  assign shiftvalin = n1145; // (signal)
  /* fppow16.vhdl:4689:8  */
  assign fixx0 = mantissa_shift_n1146; // (signal)
  /* fppow16.vhdl:4691:8  */
  assign ufixx = n1151; // (signal)
  /* fppow16.vhdl:4693:8  */
  assign expy = exp_helper_n1153; // (signal)
  /* fppow16.vhdl:4695:8  */
  assign k = exp_helper_n1154; // (signal)
  /* fppow16.vhdl:4695:11  */
  assign k_d1 = n1283; // (signal)
  /* fppow16.vhdl:4695:17  */
  assign k_d2 = n1284; // (signal)
  /* fppow16.vhdl:4697:8  */
  assign neednonorm = n1159; // (signal)
  /* fppow16.vhdl:4699:8  */
  assign preroundbiassig = n1163; // (signal)
  /* fppow16.vhdl:4701:8  */
  assign roundbit = n1168; // (signal)
  /* fppow16.vhdl:4703:8  */
  assign roundnormaddend = n1174; // (signal)
  /* fppow16.vhdl:4705:8  */
  assign roundedexpsigres = roundedexpsigoperandadder_n1176; // (signal)
  /* fppow16.vhdl:4707:8  */
  assign roundedexpsig = n1181; // (signal)
  /* fppow16.vhdl:4709:8  */
  assign ofl1 = n1189; // (signal)
  /* fppow16.vhdl:4709:14  */
  assign ofl1_d1 = n1285; // (signal)
  /* fppow16.vhdl:4709:23  */
  assign ofl1_d2 = n1286; // (signal)
  /* fppow16.vhdl:4709:32  */
  assign ofl1_d3 = n1287; // (signal)
  /* fppow16.vhdl:4709:41  */
  assign ofl1_d4 = n1288; // (signal)
  /* fppow16.vhdl:4709:50  */
  assign ofl1_d5 = n1289; // (signal)
  /* fppow16.vhdl:4711:8  */
  assign ofl2 = n1200; // (signal)
  /* fppow16.vhdl:4713:8  */
  assign ofl3 = n1206; // (signal)
  /* fppow16.vhdl:4713:14  */
  assign ofl3_d1 = n1290; // (signal)
  /* fppow16.vhdl:4713:23  */
  assign ofl3_d2 = n1291; // (signal)
  /* fppow16.vhdl:4713:32  */
  assign ofl3_d3 = n1292; // (signal)
  /* fppow16.vhdl:4713:41  */
  assign ofl3_d4 = n1293; // (signal)
  /* fppow16.vhdl:4713:50  */
  assign ofl3_d5 = n1294; // (signal)
  /* fppow16.vhdl:4713:59  */
  assign ofl3_d6 = n1295; // (signal)
  /* fppow16.vhdl:4715:8  */
  assign ofl = n1208; // (signal)
  /* fppow16.vhdl:4717:8  */
  assign ufl1 = n1216; // (signal)
  /* fppow16.vhdl:4719:8  */
  assign ufl2 = n1221; // (signal)
  /* fppow16.vhdl:4719:14  */
  assign ufl2_d1 = n1296; // (signal)
  /* fppow16.vhdl:4719:23  */
  assign ufl2_d2 = n1297; // (signal)
  /* fppow16.vhdl:4719:32  */
  assign ufl2_d3 = n1298; // (signal)
  /* fppow16.vhdl:4719:41  */
  assign ufl2_d4 = n1299; // (signal)
  /* fppow16.vhdl:4719:50  */
  assign ufl2_d5 = n1300; // (signal)
  /* fppow16.vhdl:4719:59  */
  assign ufl2_d6 = n1301; // (signal)
  /* fppow16.vhdl:4721:8  */
  assign ufl3 = n1227; // (signal)
  /* fppow16.vhdl:4721:14  */
  assign ufl3_d1 = n1302; // (signal)
  /* fppow16.vhdl:4721:23  */
  assign ufl3_d2 = n1303; // (signal)
  /* fppow16.vhdl:4721:32  */
  assign ufl3_d3 = n1304; // (signal)
  /* fppow16.vhdl:4721:41  */
  assign ufl3_d4 = n1305; // (signal)
  /* fppow16.vhdl:4721:50  */
  assign ufl3_d5 = n1306; // (signal)
  /* fppow16.vhdl:4723:8  */
  assign ufl = n1229; // (signal)
  /* fppow16.vhdl:4725:8  */
  assign rexn = n1233; // (signal)
  /* fppow16.vhdl:4801:13  */
  assign n1127 = x[25:24]; // extract
  /* fppow16.vhdl:4802:14  */
  assign n1128 = x[23]; // extract
  /* fppow16.vhdl:4803:18  */
  assign n1129 = x[22:18]; // extract
  /* fppow16.vhdl:4804:23  */
  assign n1130 = x[17:0]; // extract
  /* fppow16.vhdl:4806:22  */
  assign n1133 = {2'b00, xexpfield_d1};
  /* fppow16.vhdl:4806:38  */
  assign n1134 = n1133 - e0_d13;
  /* fppow16.vhdl:4808:31  */
  assign n1135 = shiftval[6]; // extract
  /* fppow16.vhdl:4810:15  */
  assign n1137 = {1'b1, xfrac};
  /* fppow16.vhdl:4813:29  */
  assign n1139 = shiftval[6]; // extract
  /* fppow16.vhdl:4813:17  */
  assign n1140 = ~n1139;
  /* fppow16.vhdl:4813:49  */
  assign n1141 = shiftval[5:0]; // extract
  /* fppow16.vhdl:4813:63  */
  assign n1142 = $unsigned(n1141) > $unsigned(maxshift_d13);
  /* fppow16.vhdl:4813:36  */
  assign n1143 = n1142 ? n1140 : 1'b0;
  /* fppow16.vhdl:4814:26  */
  assign n1145 = shiftval[4:0]; // extract
  /* fppow16.vhdl:4815:4  */
  leftshifter19_by_max_16_freq500_uid68 mantissa_shift (
    .clk(clk),
    .x(mxu),
    .s(shiftvalin),
    .r(mantissa_shift_n1146));
  /* fppow16.vhdl:4820:28  */
  assign n1149 = fixx0[34:18]; // extract
  /* fppow16.vhdl:4820:67  */
  assign n1150 = ~resultwillbeone_d1;
  /* fppow16.vhdl:4820:44  */
  assign n1151 = n1150 ? n1149 : 17'b00000000000000000;
  /* fppow16.vhdl:4821:4  */
  exp_5_10_freq500_uid70 exp_helper (
    .clk(clk),
    .ufixx_i(ufixx),
    .xsign(xsign),
    .expy(exp_helper_n1153),
    .k(exp_helper_n1154));
  /* fppow16.vhdl:4827:22  */
  assign n1159 = expy[13]; // extract
  /* fppow16.vhdl:4829:62  */
  assign n1160 = expy[12:3]; // extract
  /* fppow16.vhdl:4829:56  */
  assign n1162 = {7'b0001111, n1160};
  /* fppow16.vhdl:4829:76  */
  assign n1163 = neednonorm ? n1162 : n1166;
  /* fppow16.vhdl:4830:51  */
  assign n1164 = expy[11:2]; // extract
  /* fppow16.vhdl:4830:45  */
  assign n1166 = {7'b0001110, n1164};
  /* fppow16.vhdl:4831:20  */
  assign n1167 = expy[2]; // extract
  /* fppow16.vhdl:4831:25  */
  assign n1168 = neednonorm ? n1167 : n1169;
  /* fppow16.vhdl:4831:59  */
  assign n1169 = expy[1]; // extract
  /* fppow16.vhdl:4832:27  */
  assign n1170 = k_d2[5]; // extract
  /* fppow16.vhdl:4832:31  */
  assign n1171 = {n1170, k_d2};
  /* fppow16.vhdl:4832:38  */
  assign n1173 = {n1171, 9'b000000000};
  /* fppow16.vhdl:4832:60  */
  assign n1174 = {n1173, roundbit};
  /* fppow16.vhdl:4833:4  */
  intadder_17_freq500_uid111 roundedexpsigoperandadder (
    .clk(clk),
    .x(preroundbiassig),
    .y(roundnormaddend),
    .cin(n1175),
    .r(roundedexpsigoperandadder_n1176));
  /* fppow16.vhdl:4839:50  */
  assign n1180 = xexn_d6 == 2'b01;
  /* fppow16.vhdl:4839:38  */
  assign n1181 = n1180 ? roundedexpsigres : 17'b00011110000000000;
  /* fppow16.vhdl:4840:12  */
  assign n1183 = ~xsign_d1;
  /* fppow16.vhdl:4840:25  */
  assign n1184 = n1183 & overflow0;
  /* fppow16.vhdl:4840:55  */
  assign n1185 = xexn_d1[1]; // extract
  /* fppow16.vhdl:4840:44  */
  assign n1186 = ~n1185;
  /* fppow16.vhdl:4840:70  */
  assign n1187 = xexn_d1[0]; // extract
  /* fppow16.vhdl:4840:59  */
  assign n1188 = n1186 & n1187;
  /* fppow16.vhdl:4840:39  */
  assign n1189 = n1184 & n1188;
  /* fppow16.vhdl:4841:12  */
  assign n1190 = ~xsign_d6;
  /* fppow16.vhdl:4841:43  */
  assign n1191 = roundedexpsig[15]; // extract
  /* fppow16.vhdl:4841:72  */
  assign n1192 = roundedexpsig[16]; // extract
  /* fppow16.vhdl:4841:55  */
  assign n1193 = ~n1192;
  /* fppow16.vhdl:4841:51  */
  assign n1194 = n1191 & n1193;
  /* fppow16.vhdl:4841:25  */
  assign n1195 = n1190 & n1194;
  /* fppow16.vhdl:4841:99  */
  assign n1196 = xexn_d6[1]; // extract
  /* fppow16.vhdl:4841:88  */
  assign n1197 = ~n1196;
  /* fppow16.vhdl:4841:114  */
  assign n1198 = xexn_d6[0]; // extract
  /* fppow16.vhdl:4841:103  */
  assign n1199 = n1197 & n1198;
  /* fppow16.vhdl:4841:83  */
  assign n1200 = n1195 & n1199;
  /* fppow16.vhdl:4842:12  */
  assign n1201 = ~xsign;
  /* fppow16.vhdl:4842:30  */
  assign n1202 = xexn[1]; // extract
  /* fppow16.vhdl:4842:22  */
  assign n1203 = n1201 & n1202;
  /* fppow16.vhdl:4842:46  */
  assign n1204 = xexn[0]; // extract
  /* fppow16.vhdl:4842:38  */
  assign n1205 = ~n1204;
  /* fppow16.vhdl:4842:34  */
  assign n1206 = n1203 & n1205;
  /* fppow16.vhdl:4843:19  */
  assign n1207 = ofl1_d5 | ofl2;
  /* fppow16.vhdl:4843:27  */
  assign n1208 = n1207 | ofl3_d6;
  /* fppow16.vhdl:4844:26  */
  assign n1209 = roundedexpsig[15]; // extract
  /* fppow16.vhdl:4844:51  */
  assign n1210 = roundedexpsig[16]; // extract
  /* fppow16.vhdl:4844:34  */
  assign n1211 = n1209 & n1210;
  /* fppow16.vhdl:4844:79  */
  assign n1212 = xexn_d6[1]; // extract
  /* fppow16.vhdl:4844:68  */
  assign n1213 = ~n1212;
  /* fppow16.vhdl:4844:94  */
  assign n1214 = xexn_d6[0]; // extract
  /* fppow16.vhdl:4844:83  */
  assign n1215 = n1213 & n1214;
  /* fppow16.vhdl:4844:63  */
  assign n1216 = n1211 & n1215;
  /* fppow16.vhdl:4845:26  */
  assign n1217 = xexn[1]; // extract
  /* fppow16.vhdl:4845:18  */
  assign n1218 = xsign & n1217;
  /* fppow16.vhdl:4845:42  */
  assign n1219 = xexn[0]; // extract
  /* fppow16.vhdl:4845:34  */
  assign n1220 = ~n1219;
  /* fppow16.vhdl:4845:30  */
  assign n1221 = n1218 & n1220;
  /* fppow16.vhdl:4846:21  */
  assign n1222 = xsign_d1 & overflow0;
  /* fppow16.vhdl:4846:52  */
  assign n1223 = xexn_d1[1]; // extract
  /* fppow16.vhdl:4846:41  */
  assign n1224 = ~n1223;
  /* fppow16.vhdl:4846:67  */
  assign n1225 = xexn_d1[0]; // extract
  /* fppow16.vhdl:4846:56  */
  assign n1226 = n1224 & n1225;
  /* fppow16.vhdl:4846:36  */
  assign n1227 = n1222 & n1226;
  /* fppow16.vhdl:4847:16  */
  assign n1228 = ufl1 | ufl2_d6;
  /* fppow16.vhdl:4847:27  */
  assign n1229 = n1228 | ufl3_d5;
  /* fppow16.vhdl:4848:30  */
  assign n1232 = xexn_d6 == 2'b11;
  /* fppow16.vhdl:4848:17  */
  assign n1233 = n1232 ? 2'b11 : n1235;
  /* fppow16.vhdl:4849:7  */
  assign n1235 = ofl ? 2'b10 : n1237;
  /* fppow16.vhdl:4850:7  */
  assign n1237 = ufl ? 2'b00 : 2'b01;
  /* fppow16.vhdl:4852:14  */
  assign n1240 = {rexn, 1'b0};
  /* fppow16.vhdl:4852:35  */
  assign n1241 = roundedexpsig[14:0]; // extract
  /* fppow16.vhdl:4852:20  */
  assign n1242 = {n1240, n1241};
  /* fppow16.vhdl:4734:10  */
  always @(posedge clk)
    n1243 <= xexn;
  /* fppow16.vhdl:4734:10  */
  always @(posedge clk)
    n1244 <= xexn_d1;
  /* fppow16.vhdl:4734:10  */
  always @(posedge clk)
    n1245 <= xexn_d2;
  /* fppow16.vhdl:4734:10  */
  always @(posedge clk)
    n1246 <= xexn_d3;
  /* fppow16.vhdl:4734:10  */
  always @(posedge clk)
    n1247 <= xexn_d4;
  /* fppow16.vhdl:4734:10  */
  always @(posedge clk)
    n1248 <= xexn_d5;
  /* fppow16.vhdl:4734:10  */
  always @(posedge clk)
    n1249 <= xsign;
  /* fppow16.vhdl:4734:10  */
  always @(posedge clk)
    n1250 <= xsign_d1;
  /* fppow16.vhdl:4734:10  */
  always @(posedge clk)
    n1251 <= xsign_d2;
  /* fppow16.vhdl:4734:10  */
  always @(posedge clk)
    n1252 <= xsign_d3;
  /* fppow16.vhdl:4734:10  */
  always @(posedge clk)
    n1253 <= xsign_d4;
  /* fppow16.vhdl:4734:10  */
  always @(posedge clk)
    n1254 <= xsign_d5;
  /* fppow16.vhdl:4734:10  */
  always @(posedge clk)
    n1255 <= xexpfield;
  /* fppow16.vhdl:4734:10  */
  always @(posedge clk)
    n1256 <= e0;
  /* fppow16.vhdl:4734:10  */
  always @(posedge clk)
    n1257 <= e0_d1;
  /* fppow16.vhdl:4734:10  */
  always @(posedge clk)
    n1258 <= e0_d2;
  /* fppow16.vhdl:4734:10  */
  always @(posedge clk)
    n1259 <= e0_d3;
  /* fppow16.vhdl:4734:10  */
  always @(posedge clk)
    n1260 <= e0_d4;
  /* fppow16.vhdl:4734:10  */
  always @(posedge clk)
    n1261 <= e0_d5;
  /* fppow16.vhdl:4734:10  */
  always @(posedge clk)
    n1262 <= e0_d6;
  /* fppow16.vhdl:4734:10  */
  always @(posedge clk)
    n1263 <= e0_d7;
  /* fppow16.vhdl:4734:10  */
  always @(posedge clk)
    n1264 <= e0_d8;
  /* fppow16.vhdl:4734:10  */
  always @(posedge clk)
    n1265 <= e0_d9;
  /* fppow16.vhdl:4734:10  */
  always @(posedge clk)
    n1266 <= e0_d10;
  /* fppow16.vhdl:4734:10  */
  always @(posedge clk)
    n1267 <= e0_d11;
  /* fppow16.vhdl:4734:10  */
  always @(posedge clk)
    n1268 <= e0_d12;
  /* fppow16.vhdl:4734:10  */
  always @(posedge clk)
    n1269 <= resultwillbeone;
  /* fppow16.vhdl:4734:10  */
  always @(posedge clk)
    n1270 <= maxshift;
  /* fppow16.vhdl:4734:10  */
  always @(posedge clk)
    n1271 <= maxshift_d1;
  /* fppow16.vhdl:4734:10  */
  always @(posedge clk)
    n1272 <= maxshift_d2;
  /* fppow16.vhdl:4734:10  */
  always @(posedge clk)
    n1273 <= maxshift_d3;
  /* fppow16.vhdl:4734:10  */
  always @(posedge clk)
    n1274 <= maxshift_d4;
  /* fppow16.vhdl:4734:10  */
  always @(posedge clk)
    n1275 <= maxshift_d5;
  /* fppow16.vhdl:4734:10  */
  always @(posedge clk)
    n1276 <= maxshift_d6;
  /* fppow16.vhdl:4734:10  */
  always @(posedge clk)
    n1277 <= maxshift_d7;
  /* fppow16.vhdl:4734:10  */
  always @(posedge clk)
    n1278 <= maxshift_d8;
  /* fppow16.vhdl:4734:10  */
  always @(posedge clk)
    n1279 <= maxshift_d9;
  /* fppow16.vhdl:4734:10  */
  always @(posedge clk)
    n1280 <= maxshift_d10;
  /* fppow16.vhdl:4734:10  */
  always @(posedge clk)
    n1281 <= maxshift_d11;
  /* fppow16.vhdl:4734:10  */
  always @(posedge clk)
    n1282 <= maxshift_d12;
  /* fppow16.vhdl:4734:10  */
  always @(posedge clk)
    n1283 <= k;
  /* fppow16.vhdl:4734:10  */
  always @(posedge clk)
    n1284 <= k_d1;
  /* fppow16.vhdl:4734:10  */
  always @(posedge clk)
    n1285 <= ofl1;
  /* fppow16.vhdl:4734:10  */
  always @(posedge clk)
    n1286 <= ofl1_d1;
  /* fppow16.vhdl:4734:10  */
  always @(posedge clk)
    n1287 <= ofl1_d2;
  /* fppow16.vhdl:4734:10  */
  always @(posedge clk)
    n1288 <= ofl1_d3;
  /* fppow16.vhdl:4734:10  */
  always @(posedge clk)
    n1289 <= ofl1_d4;
  /* fppow16.vhdl:4734:10  */
  always @(posedge clk)
    n1290 <= ofl3;
  /* fppow16.vhdl:4734:10  */
  always @(posedge clk)
    n1291 <= ofl3_d1;
  /* fppow16.vhdl:4734:10  */
  always @(posedge clk)
    n1292 <= ofl3_d2;
  /* fppow16.vhdl:4734:10  */
  always @(posedge clk)
    n1293 <= ofl3_d3;
  /* fppow16.vhdl:4734:10  */
  always @(posedge clk)
    n1294 <= ofl3_d4;
  /* fppow16.vhdl:4734:10  */
  always @(posedge clk)
    n1295 <= ofl3_d5;
  /* fppow16.vhdl:4734:10  */
  always @(posedge clk)
    n1296 <= ufl2;
  /* fppow16.vhdl:4734:10  */
  always @(posedge clk)
    n1297 <= ufl2_d1;
  /* fppow16.vhdl:4734:10  */
  always @(posedge clk)
    n1298 <= ufl2_d2;
  /* fppow16.vhdl:4734:10  */
  always @(posedge clk)
    n1299 <= ufl2_d3;
  /* fppow16.vhdl:4734:10  */
  always @(posedge clk)
    n1300 <= ufl2_d4;
  /* fppow16.vhdl:4734:10  */
  always @(posedge clk)
    n1301 <= ufl2_d5;
  /* fppow16.vhdl:4734:10  */
  always @(posedge clk)
    n1302 <= ufl3;
  /* fppow16.vhdl:4734:10  */
  always @(posedge clk)
    n1303 <= ufl3_d1;
  /* fppow16.vhdl:4734:10  */
  always @(posedge clk)
    n1304 <= ufl3_d2;
  /* fppow16.vhdl:4734:10  */
  always @(posedge clk)
    n1305 <= ufl3_d3;
  /* fppow16.vhdl:4734:10  */
  always @(posedge clk)
    n1306 <= ufl3_d4;
endmodule

module fpmult_5_17_uid57_freq500_uid58
  (input  clk,
   input  [24:0] x,
   input  [17:0] y,
   output [25:0] r);
  wire sign;
  wire sign_d1;
  wire sign_d2;
  wire [4:0] expx;
  wire [4:0] expx_d1;
  wire [4:0] expy;
  wire [4:0] expy_d1;
  wire [4:0] expy_d2;
  wire [4:0] expy_d3;
  wire [4:0] expy_d4;
  wire [4:0] expy_d5;
  wire [4:0] expy_d6;
  wire [4:0] expy_d7;
  wire [4:0] expy_d8;
  wire [4:0] expy_d9;
  wire [4:0] expy_d10;
  wire [4:0] expy_d11;
  wire [6:0] expsumpresub;
  wire [6:0] bias;
  wire [6:0] bias_d1;
  wire [6:0] bias_d2;
  wire [6:0] bias_d3;
  wire [6:0] bias_d4;
  wire [6:0] bias_d5;
  wire [6:0] bias_d6;
  wire [6:0] bias_d7;
  wire [6:0] bias_d8;
  wire [6:0] bias_d9;
  wire [6:0] bias_d10;
  wire [6:0] bias_d11;
  wire [6:0] expsum;
  wire [17:0] sigx;
  wire [10:0] sigy;
  wire [20:0] sigprod;
  wire [3:0] excsel;
  wire [1:0] exc;
  wire [1:0] exc_d1;
  wire [1:0] exc_d2;
  wire norm;
  wire norm_d1;
  wire [6:0] exppostnorm;
  wire [20:0] sigprodext;
  wire [20:0] sigprodext_d1;
  wire [24:0] expsig;
  wire round;
  wire [24:0] expsigpostround;
  wire [1:0] excpostnorm;
  wire [1:0] finalexc;
  wire [17:0] y_d1;
  wire [17:0] y_d2;
  wire [17:0] y_d3;
  wire [17:0] y_d4;
  wire [17:0] y_d5;
  wire [17:0] y_d6;
  wire [17:0] y_d7;
  wire [17:0] y_d8;
  wire [17:0] y_d9;
  wire [17:0] y_d10;
  wire n925;
  wire n926;
  wire n927;
  wire [4:0] n928;
  wire [4:0] n929;
  wire [6:0] n931;
  wire [6:0] n933;
  wire [6:0] n934;
  wire [6:0] n936;
  wire [16:0] n937;
  wire [17:0] n939;
  wire [9:0] n940;
  wire [10:0] n942;
  wire [20:0] significandmultiplication_n943;
  wire [1:0] n946;
  wire [1:0] n947;
  wire [3:0] n948;
  wire n951;
  wire n953;
  wire n954;
  wire n956;
  wire n957;
  wire n960;
  wire n963;
  wire n965;
  wire n966;
  wire n968;
  wire n969;
  wire [2:0] n971;
  reg [1:0] n972;
  wire n973;
  wire [6:0] n975;
  wire [6:0] n976;
  wire [19:0] n977;
  wire [20:0] n979;
  wire [20:0] n980;
  wire [18:0] n981;
  wire [20:0] n983;
  wire [17:0] n984;
  wire [24:0] n985;
  localparam [24:0] n987 = 25'b0000000000000000000000000;
  wire [24:0] roundingadder_n988;
  wire [1:0] n991;
  wire n994;
  wire n997;
  wire n1000;
  wire n1002;
  wire n1003;
  wire [2:0] n1005;
  reg [1:0] n1006;
  wire n1008;
  wire n1010;
  wire n1011;
  wire n1013;
  wire n1014;
  reg [1:0] n1015;
  wire [2:0] n1016;
  wire [22:0] n1017;
  wire [25:0] n1018;
  reg n1019;
  reg n1020;
  reg [4:0] n1021;
  reg [4:0] n1022;
  reg [4:0] n1023;
  reg [4:0] n1024;
  reg [4:0] n1025;
  reg [4:0] n1026;
  reg [4:0] n1027;
  reg [4:0] n1028;
  reg [4:0] n1029;
  reg [4:0] n1030;
  reg [4:0] n1031;
  reg [4:0] n1032;
  reg [6:0] n1033;
  reg [6:0] n1034;
  reg [6:0] n1035;
  reg [6:0] n1036;
  reg [6:0] n1037;
  reg [6:0] n1038;
  reg [6:0] n1039;
  reg [6:0] n1040;
  reg [6:0] n1041;
  reg [6:0] n1042;
  reg [6:0] n1043;
  reg [1:0] n1044;
  reg [1:0] n1045;
  reg n1046;
  reg [20:0] n1047;
  reg [17:0] n1048;
  reg [17:0] n1049;
  reg [17:0] n1050;
  reg [17:0] n1051;
  reg [17:0] n1052;
  reg [17:0] n1053;
  reg [17:0] n1054;
  reg [17:0] n1055;
  reg [17:0] n1056;
  reg [17:0] n1057;
  assign r = n1018; //(module output)
  /* fppow16.vhdl:3559:8  */
  assign sign = n927; // (signal)
  /* fppow16.vhdl:3559:14  */
  assign sign_d1 = n1019; // (signal)
  /* fppow16.vhdl:3559:23  */
  assign sign_d2 = n1020; // (signal)
  /* fppow16.vhdl:3561:8  */
  assign expx = n928; // (signal)
  /* fppow16.vhdl:3561:14  */
  assign expx_d1 = n1021; // (signal)
  /* fppow16.vhdl:3563:8  */
  assign expy = n929; // (signal)
  /* fppow16.vhdl:3563:14  */
  assign expy_d1 = n1022; // (signal)
  /* fppow16.vhdl:3563:23  */
  assign expy_d2 = n1023; // (signal)
  /* fppow16.vhdl:3563:32  */
  assign expy_d3 = n1024; // (signal)
  /* fppow16.vhdl:3563:41  */
  assign expy_d4 = n1025; // (signal)
  /* fppow16.vhdl:3563:50  */
  assign expy_d5 = n1026; // (signal)
  /* fppow16.vhdl:3563:59  */
  assign expy_d6 = n1027; // (signal)
  /* fppow16.vhdl:3563:68  */
  assign expy_d7 = n1028; // (signal)
  /* fppow16.vhdl:3563:77  */
  assign expy_d8 = n1029; // (signal)
  /* fppow16.vhdl:3563:86  */
  assign expy_d9 = n1030; // (signal)
  /* fppow16.vhdl:3563:95  */
  assign expy_d10 = n1031; // (signal)
  /* fppow16.vhdl:3563:105  */
  assign expy_d11 = n1032; // (signal)
  /* fppow16.vhdl:3565:8  */
  assign expsumpresub = n934; // (signal)
  /* fppow16.vhdl:3567:8  */
  assign bias = 7'b0001111; // (signal)
  /* fppow16.vhdl:3567:14  */
  assign bias_d1 = n1033; // (signal)
  /* fppow16.vhdl:3567:23  */
  assign bias_d2 = n1034; // (signal)
  /* fppow16.vhdl:3567:32  */
  assign bias_d3 = n1035; // (signal)
  /* fppow16.vhdl:3567:41  */
  assign bias_d4 = n1036; // (signal)
  /* fppow16.vhdl:3567:50  */
  assign bias_d5 = n1037; // (signal)
  /* fppow16.vhdl:3567:59  */
  assign bias_d6 = n1038; // (signal)
  /* fppow16.vhdl:3567:68  */
  assign bias_d7 = n1039; // (signal)
  /* fppow16.vhdl:3567:77  */
  assign bias_d8 = n1040; // (signal)
  /* fppow16.vhdl:3567:86  */
  assign bias_d9 = n1041; // (signal)
  /* fppow16.vhdl:3567:95  */
  assign bias_d10 = n1042; // (signal)
  /* fppow16.vhdl:3567:105  */
  assign bias_d11 = n1043; // (signal)
  /* fppow16.vhdl:3569:8  */
  assign expsum = n936; // (signal)
  /* fppow16.vhdl:3571:8  */
  assign sigx = n939; // (signal)
  /* fppow16.vhdl:3573:8  */
  assign sigy = n942; // (signal)
  /* fppow16.vhdl:3575:8  */
  assign sigprod = significandmultiplication_n943; // (signal)
  /* fppow16.vhdl:3577:8  */
  assign excsel = n948; // (signal)
  /* fppow16.vhdl:3579:8  */
  assign exc = n972; // (signal)
  /* fppow16.vhdl:3579:13  */
  assign exc_d1 = n1044; // (signal)
  /* fppow16.vhdl:3579:21  */
  assign exc_d2 = n1045; // (signal)
  /* fppow16.vhdl:3581:8  */
  assign norm = n973; // (signal)
  /* fppow16.vhdl:3581:14  */
  assign norm_d1 = n1046; // (signal)
  /* fppow16.vhdl:3583:8  */
  assign exppostnorm = n976; // (signal)
  /* fppow16.vhdl:3585:8  */
  assign sigprodext = n980; // (signal)
  /* fppow16.vhdl:3585:20  */
  assign sigprodext_d1 = n1047; // (signal)
  /* fppow16.vhdl:3587:8  */
  assign expsig = n985; // (signal)
  /* fppow16.vhdl:3589:8  */
  assign round = 1'b1; // (signal)
  /* fppow16.vhdl:3591:8  */
  assign expsigpostround = roundingadder_n988; // (signal)
  /* fppow16.vhdl:3593:8  */
  assign excpostnorm = n1006; // (signal)
  /* fppow16.vhdl:3595:8  */
  assign finalexc = n1015; // (signal)
  /* fppow16.vhdl:3597:8  */
  assign y_d1 = n1048; // (signal)
  /* fppow16.vhdl:3597:14  */
  assign y_d2 = n1049; // (signal)
  /* fppow16.vhdl:3597:20  */
  assign y_d3 = n1050; // (signal)
  /* fppow16.vhdl:3597:26  */
  assign y_d4 = n1051; // (signal)
  /* fppow16.vhdl:3597:32  */
  assign y_d5 = n1052; // (signal)
  /* fppow16.vhdl:3597:38  */
  assign y_d6 = n1053; // (signal)
  /* fppow16.vhdl:3597:44  */
  assign y_d7 = n1054; // (signal)
  /* fppow16.vhdl:3597:50  */
  assign y_d8 = n1055; // (signal)
  /* fppow16.vhdl:3597:56  */
  assign y_d9 = n1056; // (signal)
  /* fppow16.vhdl:3597:62  */
  assign y_d10 = n1057; // (signal)
  /* fppow16.vhdl:3644:13  */
  assign n925 = x[22]; // extract
  /* fppow16.vhdl:3644:27  */
  assign n926 = y_d10[15]; // extract
  /* fppow16.vhdl:3644:18  */
  assign n927 = n925 ^ n926;
  /* fppow16.vhdl:3645:13  */
  assign n928 = x[21:17]; // extract
  /* fppow16.vhdl:3646:13  */
  assign n929 = y[14:10]; // extract
  /* fppow16.vhdl:3647:26  */
  assign n931 = {2'b00, expx_d1};
  /* fppow16.vhdl:3647:45  */
  assign n933 = {2'b00, expy_d11};
  /* fppow16.vhdl:3647:37  */
  assign n934 = n931 + n933;
  /* fppow16.vhdl:3649:27  */
  assign n936 = expsumpresub - bias_d11;
  /* fppow16.vhdl:3650:19  */
  assign n937 = x[16:0]; // extract
  /* fppow16.vhdl:3650:16  */
  assign n939 = {1'b1, n937};
  /* fppow16.vhdl:3651:19  */
  assign n940 = y[9:0]; // extract
  /* fppow16.vhdl:3651:16  */
  assign n942 = {1'b1, n940};
  /* fppow16.vhdl:3652:4  */
  intmultiplier_18x11_21_freq500_uid60 significandmultiplication (
    .clk(clk),
    .x(sigx),
    .y(sigy),
    .r(significandmultiplication_n943));
  /* fppow16.vhdl:3657:15  */
  assign n946 = x[24:23]; // extract
  /* fppow16.vhdl:3657:37  */
  assign n947 = y_d10[17:16]; // extract
  /* fppow16.vhdl:3657:30  */
  assign n948 = {n946, n947};
  /* fppow16.vhdl:3659:16  */
  assign n951 = excsel == 4'b0000;
  /* fppow16.vhdl:3659:29  */
  assign n953 = excsel == 4'b0001;
  /* fppow16.vhdl:3659:29  */
  assign n954 = n951 | n953;
  /* fppow16.vhdl:3659:38  */
  assign n956 = excsel == 4'b0100;
  /* fppow16.vhdl:3659:38  */
  assign n957 = n954 | n956;
  /* fppow16.vhdl:3660:16  */
  assign n960 = excsel == 4'b0101;
  /* fppow16.vhdl:3661:16  */
  assign n963 = excsel == 4'b0110;
  /* fppow16.vhdl:3661:28  */
  assign n965 = excsel == 4'b1001;
  /* fppow16.vhdl:3661:28  */
  assign n966 = n963 | n965;
  /* fppow16.vhdl:3661:37  */
  assign n968 = excsel == 4'b1010;
  /* fppow16.vhdl:3661:37  */
  assign n969 = n966 | n968;
  assign n971 = {n969, n960, n957};
  /* fppow16.vhdl:3658:4  */
  always @*
    case (n971)
      3'b100: n972 = 2'b10;
      3'b010: n972 = 2'b01;
      3'b001: n972 = 2'b00;
      default: n972 = 2'b11;
    endcase
  /* fppow16.vhdl:3663:19  */
  assign n973 = sigprod[20]; // extract
  /* fppow16.vhdl:3665:38  */
  assign n975 = {6'b000000, norm_d1};
  /* fppow16.vhdl:3665:26  */
  assign n976 = expsum + n975;
  /* fppow16.vhdl:3667:25  */
  assign n977 = sigprod[19:0]; // extract
  /* fppow16.vhdl:3667:39  */
  assign n979 = {n977, 1'b0};
  /* fppow16.vhdl:3667:45  */
  assign n980 = norm ? n979 : n983;
  /* fppow16.vhdl:3668:33  */
  assign n981 = sigprod[18:0]; // extract
  /* fppow16.vhdl:3668:47  */
  assign n983 = {n981, 2'b00};
  /* fppow16.vhdl:3669:41  */
  assign n984 = sigprodext_d1[20:3]; // extract
  /* fppow16.vhdl:3669:26  */
  assign n985 = {exppostnorm, n984};
  /* fppow16.vhdl:3671:4  */
  intadder_25_freq500_uid64 roundingadder (
    .clk(clk),
    .x(expsig),
    .y(n987),
    .cin(round),
    .r(roundingadder_n988));
  /* fppow16.vhdl:3677:24  */
  assign n991 = expsigpostround[24:23]; // extract
  /* fppow16.vhdl:3678:26  */
  assign n994 = n991 == 2'b00;
  /* fppow16.vhdl:3679:49  */
  assign n997 = n991 == 2'b01;
  /* fppow16.vhdl:3680:49  */
  assign n1000 = n991 == 2'b11;
  /* fppow16.vhdl:3680:58  */
  assign n1002 = n991 == 2'b10;
  /* fppow16.vhdl:3680:58  */
  assign n1003 = n1000 | n1002;
  assign n1005 = {n1003, n997, n994};
  /* fppow16.vhdl:3677:4  */
  always @*
    case (n1005)
      3'b100: n1006 = 2'b00;
      3'b010: n1006 = 2'b10;
      3'b001: n1006 = 2'b01;
      default: n1006 = 2'b11;
    endcase
  /* fppow16.vhdl:3683:23  */
  assign n1008 = exc_d2 == 2'b11;
  /* fppow16.vhdl:3683:33  */
  assign n1010 = exc_d2 == 2'b10;
  /* fppow16.vhdl:3683:33  */
  assign n1011 = n1008 | n1010;
  /* fppow16.vhdl:3683:38  */
  assign n1013 = exc_d2 == 2'b00;
  /* fppow16.vhdl:3683:38  */
  assign n1014 = n1011 | n1013;
  /* fppow16.vhdl:3682:4  */
  always @*
    case (n1014)
      1'b1: n1015 = exc_d2;
      default: n1015 = excpostnorm;
    endcase
  /* fppow16.vhdl:3685:18  */
  assign n1016 = {finalexc, sign_d2};
  /* fppow16.vhdl:3685:45  */
  assign n1017 = expsigpostround[22:0]; // extract
  /* fppow16.vhdl:3685:28  */
  assign n1018 = {n1016, n1017};
  /* fppow16.vhdl:3602:10  */
  always @(posedge clk)
    n1019 <= sign;
  /* fppow16.vhdl:3602:10  */
  always @(posedge clk)
    n1020 <= sign_d1;
  /* fppow16.vhdl:3602:10  */
  always @(posedge clk)
    n1021 <= expx;
  /* fppow16.vhdl:3602:10  */
  always @(posedge clk)
    n1022 <= expy;
  /* fppow16.vhdl:3602:10  */
  always @(posedge clk)
    n1023 <= expy_d1;
  /* fppow16.vhdl:3602:10  */
  always @(posedge clk)
    n1024 <= expy_d2;
  /* fppow16.vhdl:3602:10  */
  always @(posedge clk)
    n1025 <= expy_d3;
  /* fppow16.vhdl:3602:10  */
  always @(posedge clk)
    n1026 <= expy_d4;
  /* fppow16.vhdl:3602:10  */
  always @(posedge clk)
    n1027 <= expy_d5;
  /* fppow16.vhdl:3602:10  */
  always @(posedge clk)
    n1028 <= expy_d6;
  /* fppow16.vhdl:3602:10  */
  always @(posedge clk)
    n1029 <= expy_d7;
  /* fppow16.vhdl:3602:10  */
  always @(posedge clk)
    n1030 <= expy_d8;
  /* fppow16.vhdl:3602:10  */
  always @(posedge clk)
    n1031 <= expy_d9;
  /* fppow16.vhdl:3602:10  */
  always @(posedge clk)
    n1032 <= expy_d10;
  /* fppow16.vhdl:3602:10  */
  always @(posedge clk)
    n1033 <= bias;
  /* fppow16.vhdl:3602:10  */
  always @(posedge clk)
    n1034 <= bias_d1;
  /* fppow16.vhdl:3602:10  */
  always @(posedge clk)
    n1035 <= bias_d2;
  /* fppow16.vhdl:3602:10  */
  always @(posedge clk)
    n1036 <= bias_d3;
  /* fppow16.vhdl:3602:10  */
  always @(posedge clk)
    n1037 <= bias_d4;
  /* fppow16.vhdl:3602:10  */
  always @(posedge clk)
    n1038 <= bias_d5;
  /* fppow16.vhdl:3602:10  */
  always @(posedge clk)
    n1039 <= bias_d6;
  /* fppow16.vhdl:3602:10  */
  always @(posedge clk)
    n1040 <= bias_d7;
  /* fppow16.vhdl:3602:10  */
  always @(posedge clk)
    n1041 <= bias_d8;
  /* fppow16.vhdl:3602:10  */
  always @(posedge clk)
    n1042 <= bias_d9;
  /* fppow16.vhdl:3602:10  */
  always @(posedge clk)
    n1043 <= bias_d10;
  /* fppow16.vhdl:3602:10  */
  always @(posedge clk)
    n1044 <= exc;
  /* fppow16.vhdl:3602:10  */
  always @(posedge clk)
    n1045 <= exc_d1;
  /* fppow16.vhdl:3602:10  */
  always @(posedge clk)
    n1046 <= norm;
  /* fppow16.vhdl:3602:10  */
  always @(posedge clk)
    n1047 <= sigprodext;
  /* fppow16.vhdl:3602:10  */
  always @(posedge clk)
    n1048 <= y;
  /* fppow16.vhdl:3602:10  */
  always @(posedge clk)
    n1049 <= y_d1;
  /* fppow16.vhdl:3602:10  */
  always @(posedge clk)
    n1050 <= y_d2;
  /* fppow16.vhdl:3602:10  */
  always @(posedge clk)
    n1051 <= y_d3;
  /* fppow16.vhdl:3602:10  */
  always @(posedge clk)
    n1052 <= y_d4;
  /* fppow16.vhdl:3602:10  */
  always @(posedge clk)
    n1053 <= y_d5;
  /* fppow16.vhdl:3602:10  */
  always @(posedge clk)
    n1054 <= y_d6;
  /* fppow16.vhdl:3602:10  */
  always @(posedge clk)
    n1055 <= y_d7;
  /* fppow16.vhdl:3602:10  */
  always @(posedge clk)
    n1056 <= y_d8;
  /* fppow16.vhdl:3602:10  */
  always @(posedge clk)
    n1057 <= y_d9;
endmodule

module fplogiterative_5_17_0_500_freq500_uid9
  (input  clk,
   input  [24:0] x,
   output [24:0] r);
  wire [2:0] xexnsgn;
  wire [2:0] xexnsgn_d1;
  wire [2:0] xexnsgn_d2;
  wire [2:0] xexnsgn_d3;
  wire [2:0] xexnsgn_d4;
  wire [2:0] xexnsgn_d5;
  wire [2:0] xexnsgn_d6;
  wire [2:0] xexnsgn_d7;
  wire [2:0] xexnsgn_d8;
  wire [2:0] xexnsgn_d9;
  wire [2:0] xexnsgn_d10;
  wire firstbit;
  wire [18:0] y0;
  wire [18:0] y0_d1;
  wire [16:0] y0h;
  wire sr;
  wire sr_d1;
  wire sr_d2;
  wire sr_d3;
  wire sr_d4;
  wire sr_d5;
  wire sr_d6;
  wire sr_d7;
  wire sr_d8;
  wire sr_d9;
  wire sr_d10;
  wire [9:0] absz0;
  wire [4:0] e;
  wire [4:0] abse;
  wire eeqzero;
  wire eeqzero_d1;
  wire eeqzero_d2;
  wire eeqzero_d3;
  wire eeqzero_d4;
  wire [4:0] lzo;
  wire [4:0] lzo_d1;
  wire [4:0] lzo_d2;
  wire [4:0] lzo_d3;
  wire [4:0] pfinal_s;
  wire [4:0] pfinal_s_d1;
  wire [4:0] pfinal_s_d2;
  wire [4:0] pfinal_s_d3;
  wire [5:0] shiftval;
  wire [3:0] shiftvalinl;
  wire [3:0] shiftvalinr;
  wire dorr;
  wire dorr_d1;
  wire dorr_d2;
  wire \small ;
  wire small_d1;
  wire small_d2;
  wire small_d3;
  wire small_d4;
  wire small_d5;
  wire small_d6;
  wire [19:0] small_absz0_normd_full;
  wire [9:0] small_absz0_normd;
  wire [9:0] small_absz0_normd_d1;
  wire [6:0] a0;
  wire [7:0] inva0;
  wire [7:0] inva0_d1;
  wire [7:0] inva0_copy16;
  wire [26:0] p0;
  wire [19:0] z1;
  wire [4:0] a1;
  wire [4:0] a1_d1;
  wire [14:0] b1;
  wire [19:0] zm1;
  wire [19:0] zm1_d1;
  wire [24:0] p1;
  wire [25:0] y1;
  wire [20:0] eiy1;
  wire [20:0] addxiter1;
  wire [20:0] eiypb1;
  wire [20:0] pp1;
  wire [20:0] z2;
  wire [20:0] zfinal;
  wire [20:0] zfinal_d1;
  wire [20:0] zfinal_d2;
  wire [13:0] squarerin;
  wire [27:0] z2o2_full;
  wire [27:0] z2o2_full_dummy;
  wire [10:0] z2o2_normal;
  wire [20:0] addfinallog1py;
  wire [20:0] log1p_normal;
  wire [29:0] l0;
  wire [29:0] l0_copy28;
  wire [29:0] s1;
  wire [24:0] l1;
  wire [24:0] l1_copy31;
  wire [29:0] sopx1;
  wire [29:0] s2;
  wire [29:0] almostlog;
  wire [29:0] adderlogf_normaly;
  wire [29:0] logf_normal;
  wire [25:0] abselog2;
  wire [34:0] abselog2_pad;
  wire [34:0] logf_normal_pad;
  wire [34:0] lnaddx;
  wire [34:0] lnaddy;
  wire [34:0] log_normal;
  wire [29:0] log_normal_normd;
  wire [29:0] log_normal_normd_d1;
  wire [3:0] e_normal;
  wire [13:0] z2o2_small_bs;
  wire [26:0] z2o2_small_s;
  wire [22:0] z2o2_small;
  wire [22:0] z_small;
  wire [22:0] log_smally;
  wire nsrcin;
  wire [22:0] log_small;
  wire [1:0] e0_sub;
  wire [5:0] e_small;
  wire [5:0] e_small_d1;
  wire [5:0] e_small_d2;
  wire [5:0] e_small_d3;
  wire ufl;
  wire ufl_d1;
  wire ufl_d2;
  wire ufl_d3;
  wire ufl_d4;
  wire [20:0] log_small_normd;
  wire [20:0] log_small_normd_d1;
  wire [20:0] log_small_normd_d2;
  wire [20:0] log_small_normd_d3;
  wire [20:0] log_small_normd_d4;
  wire [4:0] e0offset;
  wire [4:0] e0offset_d1;
  wire [4:0] e0offset_d2;
  wire [4:0] e0offset_d3;
  wire [4:0] e0offset_d4;
  wire [4:0] e0offset_d5;
  wire [4:0] e0offset_d6;
  wire [4:0] e0offset_d7;
  wire [4:0] e0offset_d8;
  wire [4:0] e0offset_d9;
  wire [4:0] er;
  wire [20:0] log_g;
  wire round;
  wire [21:0] frax;
  wire [21:0] fray;
  wire [21:0] efr;
  wire [2:0] rexn;
  wire [2:0] n569;
  wire n570;
  wire [16:0] n571;
  wire [17:0] n573;
  wire [18:0] n575;
  wire n576;
  wire [18:0] n577;
  wire [16:0] n578;
  wire [18:0] n580;
  wire [16:0] n581;
  wire [4:0] n583;
  wire n585;
  wire n586;
  wire n587;
  wire n588;
  wire [9:0] n589;
  wire n590;
  wire [9:0] n591;
  wire [9:0] n592;
  wire [9:0] n594;
  wire [4:0] n595;
  wire n596;
  wire [4:0] n598;
  wire [4:0] n599;
  wire [4:0] n601;
  wire [4:0] n602;
  wire n605;
  wire n606;
  wire [4:0] lzoc1_n608;
  wire [5:0] n613;
  wire [5:0] n615;
  wire [5:0] n616;
  wire [3:0] n617;
  wire [3:0] n618;
  wire n619;
  wire n620;
  wire n621;
  wire [19:0] small_lshift_n622;
  wire [9:0] n625;
  wire [6:0] n626;
  wire [7:0] inva0table_n627;
  wire [26:0] n630;
  wire [26:0] n631;
  wire [26:0] n632;
  wire [19:0] n633;
  wire [4:0] n634;
  wire [14:0] n635;
  wire [24:0] n636;
  wire [24:0] n637;
  wire [24:0] n638;
  wire [25:0] n640;
  wire [20:0] n641;
  wire n642;
  wire [20:0] n643;
  wire [19:0] n644;
  wire [20:0] n646;
  wire [15:0] n648;
  wire [20:0] n650;
  localparam n651 = 1'b0;
  wire [20:0] additer1_1_n652;
  wire [19:0] n655;
  wire [19:0] n656;
  wire [20:0] n658;
  localparam n659 = 1'b1;
  wire [20:0] additer2_1_n660;
  wire [13:0] n663;
  wire [13:0] n664;
  wire [13:0] n666;
  wire [27:0] n667;
  wire [27:0] n668;
  wire [27:0] n669;
  wire [10:0] n670;
  wire [10:0] n671;
  wire [20:0] n673;
  localparam n674 = 1'b1;
  wire [20:0] addfinallog1p_normaladder_n675;
  wire [29:0] logtable0_n678;
  wire [24:0] logtable1_n681;
  wire [29:0] n685;
  localparam n686 = 1'b0;
  wire [29:0] adders1_n687;
  wire [29:0] n691;
  localparam n692 = 1'b0;
  wire [29:0] adderlogf_normal_n693;
  wire [25:0] mullog2_n696;
  wire [34:0] n700;
  wire n701;
  wire n702;
  wire n703;
  wire n704;
  wire n705;
  wire [3:0] n706;
  wire [4:0] n707;
  wire [34:0] n708;
  wire n709;
  wire [34:0] n710;
  wire [34:0] n711;
  wire [34:0] lnadder_n712;
  wire [3:0] final_norm_n715;
  wire [29:0] final_norm_n716;
  wire [13:0] n721;
  wire [26:0] ao_rshift_n722;
  wire [13:0] n725;
  wire [22:0] n727;
  wire [22:0] n729;
  wire [22:0] n730;
  wire [22:0] n731;
  wire n732;
  wire [22:0] log_small_adder_n733;
  wire n737;
  wire [1:0] n738;
  wire [1:0] n740;
  wire n742;
  wire [1:0] n743;
  wire [5:0] n746;
  wire [5:0] n748;
  wire [5:0] n749;
  wire n750;
  wire [20:0] n751;
  wire n752;
  wire [20:0] n753;
  wire [20:0] n754;
  wire n755;
  wire [20:0] n756;
  wire [20:0] n757;
  wire [4:0] n759;
  wire [4:0] n760;
  wire [4:0] n762;
  wire [4:0] n763;
  wire [19:0] n764;
  wire [20:0] n766;
  wire [20:0] n767;
  wire [20:0] n768;
  wire n769;
  wire [16:0] n770;
  wire [21:0] n771;
  wire [21:0] n773;
  localparam n774 = 1'b0;
  wire [21:0] finalroundadder_n775;
  wire n779;
  wire n780;
  wire n781;
  wire n782;
  wire n783;
  wire n784;
  wire n785;
  wire n786;
  wire n787;
  wire [2:0] n788;
  wire [1:0] n790;
  wire n792;
  wire [2:0] n793;
  wire [1:0] n795;
  wire n797;
  wire [2:0] n798;
  wire [2:0] n800;
  wire n801;
  wire n802;
  wire n803;
  wire n804;
  wire n805;
  wire n806;
  wire n807;
  wire n808;
  wire n809;
  wire n810;
  wire [2:0] n811;
  wire [2:0] n813;
  wire [24:0] n814;
  reg [2:0] n815;
  reg [2:0] n816;
  reg [2:0] n817;
  reg [2:0] n818;
  reg [2:0] n819;
  reg [2:0] n820;
  reg [2:0] n821;
  reg [2:0] n822;
  reg [2:0] n823;
  reg [2:0] n824;
  reg [18:0] n825;
  reg n826;
  reg n827;
  reg n828;
  reg n829;
  reg n830;
  reg n831;
  reg n832;
  reg n833;
  reg n834;
  reg n835;
  reg n836;
  reg n837;
  reg n838;
  reg n839;
  reg [4:0] n840;
  reg [4:0] n841;
  reg [4:0] n842;
  reg [4:0] n843;
  reg [4:0] n844;
  reg [4:0] n845;
  reg n846;
  reg n847;
  reg n848;
  reg n849;
  reg n850;
  reg n851;
  reg n852;
  reg n853;
  reg [9:0] n854;
  reg [7:0] n855;
  reg [4:0] n856;
  reg [19:0] n857;
  reg [20:0] n858;
  reg [20:0] n859;
  reg [29:0] n860;
  reg [5:0] n861;
  reg [5:0] n862;
  reg [5:0] n863;
  reg n864;
  reg n865;
  reg n866;
  reg n867;
  reg [20:0] n868;
  reg [20:0] n869;
  reg [20:0] n870;
  reg [20:0] n871;
  reg [4:0] n872;
  reg [4:0] n873;
  reg [4:0] n874;
  reg [4:0] n875;
  reg [4:0] n876;
  reg [4:0] n877;
  reg [4:0] n878;
  reg [4:0] n879;
  reg [4:0] n880;
  assign r = n814; //(module output)
  /* fppow16.vhdl:2968:8  */
  assign xexnsgn = n569; // (signal)
  /* fppow16.vhdl:2968:17  */
  assign xexnsgn_d1 = n815; // (signal)
  /* fppow16.vhdl:2968:29  */
  assign xexnsgn_d2 = n816; // (signal)
  /* fppow16.vhdl:2968:41  */
  assign xexnsgn_d3 = n817; // (signal)
  /* fppow16.vhdl:2968:53  */
  assign xexnsgn_d4 = n818; // (signal)
  /* fppow16.vhdl:2968:65  */
  assign xexnsgn_d5 = n819; // (signal)
  /* fppow16.vhdl:2968:77  */
  assign xexnsgn_d6 = n820; // (signal)
  /* fppow16.vhdl:2968:89  */
  assign xexnsgn_d7 = n821; // (signal)
  /* fppow16.vhdl:2968:101  */
  assign xexnsgn_d8 = n822; // (signal)
  /* fppow16.vhdl:2968:113  */
  assign xexnsgn_d9 = n823; // (signal)
  /* fppow16.vhdl:2968:125  */
  assign xexnsgn_d10 = n824; // (signal)
  /* fppow16.vhdl:2970:8  */
  assign firstbit = n570; // (signal)
  /* fppow16.vhdl:2972:8  */
  assign y0 = n577; // (signal)
  /* fppow16.vhdl:2972:12  */
  assign y0_d1 = n825; // (signal)
  /* fppow16.vhdl:2974:8  */
  assign y0h = n581; // (signal)
  /* fppow16.vhdl:2976:8  */
  assign sr = n586; // (signal)
  /* fppow16.vhdl:2976:12  */
  assign sr_d1 = n826; // (signal)
  /* fppow16.vhdl:2976:19  */
  assign sr_d2 = n827; // (signal)
  /* fppow16.vhdl:2976:26  */
  assign sr_d3 = n828; // (signal)
  /* fppow16.vhdl:2976:33  */
  assign sr_d4 = n829; // (signal)
  /* fppow16.vhdl:2976:40  */
  assign sr_d5 = n830; // (signal)
  /* fppow16.vhdl:2976:47  */
  assign sr_d6 = n831; // (signal)
  /* fppow16.vhdl:2976:54  */
  assign sr_d7 = n832; // (signal)
  /* fppow16.vhdl:2976:61  */
  assign sr_d8 = n833; // (signal)
  /* fppow16.vhdl:2976:68  */
  assign sr_d9 = n834; // (signal)
  /* fppow16.vhdl:2976:75  */
  assign sr_d10 = n835; // (signal)
  /* fppow16.vhdl:2978:8  */
  assign absz0 = n591; // (signal)
  /* fppow16.vhdl:2980:8  */
  assign e = n599; // (signal)
  /* fppow16.vhdl:2982:8  */
  assign abse = n602; // (signal)
  /* fppow16.vhdl:2984:8  */
  assign eeqzero = n606; // (signal)
  /* fppow16.vhdl:2984:17  */
  assign eeqzero_d1 = n836; // (signal)
  /* fppow16.vhdl:2984:29  */
  assign eeqzero_d2 = n837; // (signal)
  /* fppow16.vhdl:2984:41  */
  assign eeqzero_d3 = n838; // (signal)
  /* fppow16.vhdl:2984:53  */
  assign eeqzero_d4 = n839; // (signal)
  /* fppow16.vhdl:2986:8  */
  assign lzo = lzoc1_n608; // (signal)
  /* fppow16.vhdl:2986:13  */
  assign lzo_d1 = n840; // (signal)
  /* fppow16.vhdl:2986:21  */
  assign lzo_d2 = n841; // (signal)
  /* fppow16.vhdl:2986:29  */
  assign lzo_d3 = n842; // (signal)
  /* fppow16.vhdl:2988:8  */
  assign pfinal_s = 5'b01001; // (signal)
  /* fppow16.vhdl:2988:18  */
  assign pfinal_s_d1 = n843; // (signal)
  /* fppow16.vhdl:2988:31  */
  assign pfinal_s_d2 = n844; // (signal)
  /* fppow16.vhdl:2988:44  */
  assign pfinal_s_d3 = n845; // (signal)
  /* fppow16.vhdl:2990:8  */
  assign shiftval = n616; // (signal)
  /* fppow16.vhdl:2992:8  */
  assign shiftvalinl = n617; // (signal)
  /* fppow16.vhdl:2994:8  */
  assign shiftvalinr = n618; // (signal)
  /* fppow16.vhdl:2996:8  */
  assign dorr = n619; // (signal)
  /* fppow16.vhdl:2996:14  */
  assign dorr_d1 = n846; // (signal)
  /* fppow16.vhdl:2996:23  */
  assign dorr_d2 = n847; // (signal)
  /* fppow16.vhdl:2998:8  */
  assign \small  = n621; // (signal)
  /* fppow16.vhdl:2998:15  */
  assign small_d1 = n848; // (signal)
  /* fppow16.vhdl:2998:25  */
  assign small_d2 = n849; // (signal)
  /* fppow16.vhdl:2998:35  */
  assign small_d3 = n850; // (signal)
  /* fppow16.vhdl:2998:45  */
  assign small_d4 = n851; // (signal)
  /* fppow16.vhdl:2998:55  */
  assign small_d5 = n852; // (signal)
  /* fppow16.vhdl:2998:65  */
  assign small_d6 = n853; // (signal)
  /* fppow16.vhdl:3000:8  */
  assign small_absz0_normd_full = small_lshift_n622; // (signal)
  /* fppow16.vhdl:3002:8  */
  assign small_absz0_normd = n625; // (signal)
  /* fppow16.vhdl:3002:27  */
  assign small_absz0_normd_d1 = n854; // (signal)
  /* fppow16.vhdl:3004:8  */
  assign a0 = n626; // (signal)
  /* fppow16.vhdl:3006:8  */
  assign inva0 = inva0_copy16; // (signal)
  /* fppow16.vhdl:3006:15  */
  assign inva0_d1 = n855; // (signal)
  /* fppow16.vhdl:3008:8  */
  assign inva0_copy16 = inva0table_n627; // (signal)
  /* fppow16.vhdl:3010:8  */
  assign p0 = n632; // (signal)
  /* fppow16.vhdl:3012:8  */
  assign z1 = n633; // (signal)
  /* fppow16.vhdl:3014:8  */
  assign a1 = n634; // (signal)
  /* fppow16.vhdl:3014:12  */
  assign a1_d1 = n856; // (signal)
  /* fppow16.vhdl:3016:8  */
  assign b1 = n635; // (signal)
  /* fppow16.vhdl:3018:8  */
  assign zm1 = z1; // (signal)
  /* fppow16.vhdl:3018:13  */
  assign zm1_d1 = n857; // (signal)
  /* fppow16.vhdl:3020:8  */
  assign p1 = n638; // (signal)
  /* fppow16.vhdl:3022:8  */
  assign y1 = n640; // (signal)
  /* fppow16.vhdl:3024:8  */
  assign eiy1 = n643; // (signal)
  /* fppow16.vhdl:3026:8  */
  assign addxiter1 = n650; // (signal)
  /* fppow16.vhdl:3028:8  */
  assign eiypb1 = additer1_1_n652; // (signal)
  /* fppow16.vhdl:3030:8  */
  assign pp1 = n658; // (signal)
  /* fppow16.vhdl:3032:8  */
  assign z2 = additer2_1_n660; // (signal)
  /* fppow16.vhdl:3034:8  */
  assign zfinal = z2; // (signal)
  /* fppow16.vhdl:3034:16  */
  assign zfinal_d1 = n858; // (signal)
  /* fppow16.vhdl:3034:27  */
  assign zfinal_d2 = n859; // (signal)
  /* fppow16.vhdl:3036:8  */
  assign squarerin = n664; // (signal)
  /* fppow16.vhdl:3038:8  */
  assign z2o2_full = n669; // (signal)
  /* fppow16.vhdl:3040:8  */
  assign z2o2_full_dummy = z2o2_full; // (signal)
  /* fppow16.vhdl:3042:8  */
  assign z2o2_normal = n670; // (signal)
  /* fppow16.vhdl:3044:8  */
  assign addfinallog1py = n673; // (signal)
  /* fppow16.vhdl:3046:8  */
  assign log1p_normal = addfinallog1p_normaladder_n675; // (signal)
  /* fppow16.vhdl:3048:8  */
  assign l0 = l0_copy28; // (signal)
  /* fppow16.vhdl:3050:8  */
  assign l0_copy28 = logtable0_n678; // (signal)
  /* fppow16.vhdl:3052:8  */
  assign s1 = l0; // (signal)
  /* fppow16.vhdl:3054:8  */
  assign l1 = l1_copy31; // (signal)
  /* fppow16.vhdl:3056:8  */
  assign l1_copy31 = logtable1_n681; // (signal)
  /* fppow16.vhdl:3058:8  */
  assign sopx1 = n685; // (signal)
  /* fppow16.vhdl:3060:8  */
  assign s2 = adders1_n687; // (signal)
  /* fppow16.vhdl:3062:8  */
  assign almostlog = s2; // (signal)
  /* fppow16.vhdl:3064:8  */
  assign adderlogf_normaly = n691; // (signal)
  /* fppow16.vhdl:3066:8  */
  assign logf_normal = adderlogf_normal_n693; // (signal)
  /* fppow16.vhdl:3068:8  */
  assign abselog2 = mullog2_n696; // (signal)
  /* fppow16.vhdl:3070:8  */
  assign abselog2_pad = n700; // (signal)
  /* fppow16.vhdl:3072:8  */
  assign logf_normal_pad = n708; // (signal)
  /* fppow16.vhdl:3074:8  */
  assign lnaddx = abselog2_pad; // (signal)
  /* fppow16.vhdl:3076:8  */
  assign lnaddy = n710; // (signal)
  /* fppow16.vhdl:3078:8  */
  assign log_normal = lnadder_n712; // (signal)
  /* fppow16.vhdl:3080:8  */
  assign log_normal_normd = final_norm_n716; // (signal)
  /* fppow16.vhdl:3080:26  */
  assign log_normal_normd_d1 = n860; // (signal)
  /* fppow16.vhdl:3082:8  */
  assign e_normal = final_norm_n715; // (signal)
  /* fppow16.vhdl:3084:8  */
  assign z2o2_small_bs = n721; // (signal)
  /* fppow16.vhdl:3086:8  */
  assign z2o2_small_s = ao_rshift_n722; // (signal)
  /* fppow16.vhdl:3088:8  */
  assign z2o2_small = n727; // (signal)
  /* fppow16.vhdl:3090:8  */
  assign z_small = n729; // (signal)
  /* fppow16.vhdl:3092:8  */
  assign log_smally = n730; // (signal)
  /* fppow16.vhdl:3094:8  */
  assign nsrcin = n732; // (signal)
  /* fppow16.vhdl:3096:8  */
  assign log_small = log_small_adder_n733; // (signal)
  /* fppow16.vhdl:3098:8  */
  assign e0_sub = n738; // (signal)
  /* fppow16.vhdl:3100:8  */
  assign e_small = n749; // (signal)
  /* fppow16.vhdl:3100:17  */
  assign e_small_d1 = n861; // (signal)
  /* fppow16.vhdl:3100:29  */
  assign e_small_d2 = n862; // (signal)
  /* fppow16.vhdl:3100:41  */
  assign e_small_d3 = n863; // (signal)
  /* fppow16.vhdl:3102:8  */
  assign ufl = n750; // (signal)
  /* fppow16.vhdl:3102:13  */
  assign ufl_d1 = n864; // (signal)
  /* fppow16.vhdl:3102:21  */
  assign ufl_d2 = n865; // (signal)
  /* fppow16.vhdl:3102:29  */
  assign ufl_d3 = n866; // (signal)
  /* fppow16.vhdl:3102:37  */
  assign ufl_d4 = n867; // (signal)
  /* fppow16.vhdl:3104:8  */
  assign log_small_normd = n753; // (signal)
  /* fppow16.vhdl:3104:25  */
  assign log_small_normd_d1 = n868; // (signal)
  /* fppow16.vhdl:3104:45  */
  assign log_small_normd_d2 = n869; // (signal)
  /* fppow16.vhdl:3104:65  */
  assign log_small_normd_d3 = n870; // (signal)
  /* fppow16.vhdl:3104:85  */
  assign log_small_normd_d4 = n871; // (signal)
  /* fppow16.vhdl:3106:8  */
  assign e0offset = 5'b10011; // (signal)
  /* fppow16.vhdl:3106:18  */
  assign e0offset_d1 = n872; // (signal)
  /* fppow16.vhdl:3106:31  */
  assign e0offset_d2 = n873; // (signal)
  /* fppow16.vhdl:3106:44  */
  assign e0offset_d3 = n874; // (signal)
  /* fppow16.vhdl:3106:57  */
  assign e0offset_d4 = n875; // (signal)
  /* fppow16.vhdl:3106:70  */
  assign e0offset_d5 = n876; // (signal)
  /* fppow16.vhdl:3106:83  */
  assign e0offset_d6 = n877; // (signal)
  /* fppow16.vhdl:3106:96  */
  assign e0offset_d7 = n878; // (signal)
  /* fppow16.vhdl:3106:109  */
  assign e0offset_d8 = n879; // (signal)
  /* fppow16.vhdl:3106:122  */
  assign e0offset_d9 = n880; // (signal)
  /* fppow16.vhdl:3108:8  */
  assign er = n760; // (signal)
  /* fppow16.vhdl:3110:8  */
  assign log_g = n767; // (signal)
  /* fppow16.vhdl:3112:8  */
  assign round = n769; // (signal)
  /* fppow16.vhdl:3114:8  */
  assign frax = n771; // (signal)
  /* fppow16.vhdl:3116:8  */
  assign fray = n773; // (signal)
  /* fppow16.vhdl:3118:8  */
  assign efr = finalroundadder_n775; // (signal)
  /* fppow16.vhdl:3120:8  */
  assign rexn = n788; // (signal)
  /* fppow16.vhdl:3201:17  */
  assign n569 = x[24:22]; // extract
  /* fppow16.vhdl:3202:18  */
  assign n570 = x[16]; // extract
  /* fppow16.vhdl:3203:17  */
  assign n571 = x[16:0]; // extract
  /* fppow16.vhdl:3203:14  */
  assign n573 = {1'b1, n571};
  /* fppow16.vhdl:3203:33  */
  assign n575 = {n573, 1'b0};
  /* fppow16.vhdl:3203:53  */
  assign n576 = ~firstbit;
  /* fppow16.vhdl:3203:39  */
  assign n577 = n576 ? n575 : n580;
  /* fppow16.vhdl:3203:72  */
  assign n578 = x[16:0]; // extract
  /* fppow16.vhdl:3203:69  */
  assign n580 = {2'b01, n578};
  /* fppow16.vhdl:3204:13  */
  assign n581 = y0[17:1]; // extract
  /* fppow16.vhdl:3206:24  */
  assign n583 = x[21:17]; // extract
  /* fppow16.vhdl:3206:44  */
  assign n585 = n583 == 5'b01111;
  /* fppow16.vhdl:3206:16  */
  assign n586 = n585 ? 1'b0 : n588;
  /* fppow16.vhdl:3207:16  */
  assign n587 = x[21]; // extract
  /* fppow16.vhdl:3207:11  */
  assign n588 = ~n587;
  /* fppow16.vhdl:3208:17  */
  assign n589 = y0[9:0]; // extract
  /* fppow16.vhdl:3208:57  */
  assign n590 = ~sr;
  /* fppow16.vhdl:3208:49  */
  assign n591 = n590 ? n589 : n594;
  /* fppow16.vhdl:3209:49  */
  assign n592 = y0[9:0]; // extract
  /* fppow16.vhdl:3209:45  */
  assign n594 = 10'b0000000000 - n592;
  /* fppow16.vhdl:3210:11  */
  assign n595 = x[21:17]; // extract
  /* fppow16.vhdl:3210:67  */
  assign n596 = ~firstbit;
  /* fppow16.vhdl:3210:64  */
  assign n598 = {4'b0111, n596};
  /* fppow16.vhdl:3210:32  */
  assign n599 = n595 - n598;
  /* fppow16.vhdl:3211:36  */
  assign n601 = 5'b00000 - e;
  /* fppow16.vhdl:3211:43  */
  assign n602 = sr ? n601 : e;
  /* fppow16.vhdl:3212:25  */
  assign n605 = e == 5'b00000;
  /* fppow16.vhdl:3212:19  */
  assign n606 = n605 ? 1'b1 : 1'b0;
  /* fppow16.vhdl:3213:4  */
  lzoc_17_freq500_uid11 lzoc1 (
    .clk(clk),
    .i(y0h),
    .ozb(firstbit),
    .o(lzoc1_n608));
  /* fppow16.vhdl:3219:21  */
  assign n613 = {1'b0, lzo};
  /* fppow16.vhdl:3219:35  */
  assign n615 = {1'b0, pfinal_s_d3};
  /* fppow16.vhdl:3219:28  */
  assign n616 = n613 - n615;
  /* fppow16.vhdl:3220:27  */
  assign n617 = shiftval[3:0]; // extract
  /* fppow16.vhdl:3221:27  */
  assign n618 = shiftval[3:0]; // extract
  /* fppow16.vhdl:3222:20  */
  assign n619 = shiftval[5]; // extract
  /* fppow16.vhdl:3223:28  */
  assign n620 = ~dorr_d1;
  /* fppow16.vhdl:3223:24  */
  assign n621 = eeqzero_d4 & n620;
  /* fppow16.vhdl:3225:4  */
  leftshifter10_by_max_10_freq500_uid13 small_lshift (
    .clk(clk),
    .x(absz0),
    .s(shiftvalinl),
    .r(small_lshift_n622));
  /* fppow16.vhdl:3230:47  */
  assign n625 = small_absz0_normd_full[9:0]; // extract
  /* fppow16.vhdl:3232:11  */
  assign n626 = x[16:10]; // extract
  /* fppow16.vhdl:3234:4  */
  inva0table_freq500_uid15 inva0table (
    .x(a0),
    .y(inva0table_n627));
  /* fppow16.vhdl:3238:19  */
  assign n630 = {19'b0, inva0_d1};  //  uext
  /* fppow16.vhdl:3238:19  */
  assign n631 = {8'b0, y0_d1};  //  uext
  /* fppow16.vhdl:3238:19  */
  assign n632 = n630 * n631; // umul
  /* fppow16.vhdl:3240:12  */
  assign n633 = p0[19:0]; // extract
  /* fppow16.vhdl:3242:12  */
  assign n634 = z1[19:15]; // extract
  /* fppow16.vhdl:3243:12  */
  assign n635 = z1[14:0]; // extract
  /* fppow16.vhdl:3245:15  */
  assign n636 = {20'b0, a1_d1};  //  uext
  /* fppow16.vhdl:3245:15  */
  assign n637 = {5'b0, zm1_d1};  //  uext
  /* fppow16.vhdl:3245:15  */
  assign n638 = n636 * n637; // umul
  /* fppow16.vhdl:3246:36  */
  assign n640 = {6'b100000, z1};
  /* fppow16.vhdl:3247:14  */
  assign n641 = y1[25:5]; // extract
  /* fppow16.vhdl:3247:36  */
  assign n642 = a1[4]; // extract
  /* fppow16.vhdl:3247:29  */
  assign n643 = n642 ? n641 : n646;
  /* fppow16.vhdl:3248:20  */
  assign n644 = y1[25:6]; // extract
  /* fppow16.vhdl:3248:16  */
  assign n646 = {1'b0, n644};
  /* fppow16.vhdl:3249:21  */
  assign n648 = {1'b0, b1};
  /* fppow16.vhdl:3249:26  */
  assign n650 = {n648, 5'b00000};
  /* fppow16.vhdl:3250:4  */
  intadder_21_freq500_uid19 additer1_1 (
    .clk(clk),
    .x(addxiter1),
    .y(eiy1),
    .cin(n651),
    .r(additer1_1_n652));
  /* fppow16.vhdl:3256:39  */
  assign n655 = p1[24:5]; // extract
  /* fppow16.vhdl:3256:33  */
  assign n656 = ~n655;
  /* fppow16.vhdl:3256:31  */
  assign n658 = {1'b1, n656};
  /* fppow16.vhdl:3257:4  */
  intadder_21_freq500_uid22 additer2_1 (
    .clk(clk),
    .x(eiypb1),
    .y(pp1),
    .cin(n659),
    .r(additer2_1_n660));
  /* fppow16.vhdl:3264:26  */
  assign n663 = zfinal_d2[20:7]; // extract
  /* fppow16.vhdl:3264:54  */
  assign n664 = dorr_d2 ? n663 : n666;
  /* fppow16.vhdl:3265:48  */
  assign n666 = {small_absz0_normd_d1, 4'b0000};
  /* fppow16.vhdl:3266:26  */
  assign n667 = {14'b0, squarerin};  //  uext
  /* fppow16.vhdl:3266:26  */
  assign n668 = {14'b0, squarerin};  //  uext
  /* fppow16.vhdl:3266:26  */
  assign n669 = n667 * n668; // umul
  /* fppow16.vhdl:3268:35  */
  assign n670 = z2o2_full_dummy[27:17]; // extract
  /* fppow16.vhdl:3269:50  */
  assign n671 = ~z2o2_normal;
  /* fppow16.vhdl:3269:48  */
  assign n673 = {10'b1111111111, n671};
  /* fppow16.vhdl:3270:4  */
  intadder_21_freq500_uid25 addfinallog1p_normaladder (
    .clk(clk),
    .x(zfinal),
    .y(addfinallog1py),
    .cin(n674),
    .r(addfinallog1p_normaladder_n675));
  /* fppow16.vhdl:3278:4  */
  logtable0_freq500_uid27 logtable0 (
    .x(a0),
    .y(logtable0_n678));
  /* fppow16.vhdl:3283:4  */
  logtable1_freq500_uid30 logtable1 (
    .x(a1),
    .y(logtable1_n681));
  /* fppow16.vhdl:3287:36  */
  assign n685 = {5'b00000, l1};
  /* fppow16.vhdl:3288:4  */
  intadder_30_freq500_uid34 adders1 (
    .clk(clk),
    .x(s1),
    .y(sopx1),
    .cin(n686),
    .r(adders1_n687));
  /* fppow16.vhdl:3295:62  */
  assign n691 = {9'b000000000, log1p_normal};
  /* fppow16.vhdl:3296:4  */
  intadder_30_freq500_uid37 adderlogf_normal (
    .clk(clk),
    .x(almostlog),
    .y(adderlogf_normaly),
    .cin(n692),
    .r(adderlogf_normal_n693));
  /* fppow16.vhdl:3302:4  */
  fixrealkcm_freq500_uid39 mullog2 (
    .clk(clk),
    .x(abse),
    .r(mullog2_n696));
  /* fppow16.vhdl:3306:31  */
  assign n700 = {abselog2, 9'b000000000};
  /* fppow16.vhdl:3307:53  */
  assign n701 = logf_normal[29]; // extract
  /* fppow16.vhdl:3307:53  */
  assign n702 = logf_normal[29]; // extract
  /* fppow16.vhdl:3307:53  */
  assign n703 = logf_normal[29]; // extract
  /* fppow16.vhdl:3307:53  */
  assign n704 = logf_normal[29]; // extract
  /* fppow16.vhdl:3307:53  */
  assign n705 = logf_normal[29]; // extract
  assign n706 = {n705, n704, n703, n702};
  assign n707 = {n706, n701};
  /* fppow16.vhdl:3307:70  */
  assign n708 = {n707, logf_normal};
  /* fppow16.vhdl:3309:40  */
  assign n709 = ~sr_d6;
  /* fppow16.vhdl:3309:30  */
  assign n710 = n709 ? logf_normal_pad : n711;
  /* fppow16.vhdl:3309:50  */
  assign n711 = ~logf_normal_pad;
  /* fppow16.vhdl:3310:4  */
  intadder_35_freq500_uid46 lnadder (
    .clk(clk),
    .x(lnaddx),
    .y(lnaddy),
    .cin(sr),
    .r(lnadder_n712));
  /* fppow16.vhdl:3316:4  */
  normalizer_z_35_30_13_freq500_uid48 final_norm (
    .clk(clk),
    .x(log_normal),
    .count(final_norm_n715),
    .r(final_norm_n716));
  /* fppow16.vhdl:3321:36  */
  assign n721 = z2o2_full_dummy[27:14]; // extract
  /* fppow16.vhdl:3322:4  */
  rightshifter14_by_max_13_freq500_uid50 ao_rshift (
    .clk(clk),
    .x(z2o2_small_bs),
    .s(shiftvalinr),
    .r(ao_rshift_n722));
  /* fppow16.vhdl:3328:61  */
  assign n725 = z2o2_small_s[26:13]; // extract
  /* fppow16.vhdl:3328:47  */
  assign n727 = {9'b000000000, n725};
  /* fppow16.vhdl:3330:33  */
  assign n729 = {small_absz0_normd, 13'b0000000000000};
  /* fppow16.vhdl:3331:29  */
  assign n730 = sr_d6 ? z2o2_small : n731;
  /* fppow16.vhdl:3331:49  */
  assign n731 = ~z2o2_small;
  /* fppow16.vhdl:3332:14  */
  assign n732 = ~sr;
  /* fppow16.vhdl:3333:4  */
  intadder_23_freq500_uid52 log_small_adder (
    .clk(clk),
    .x(z_small),
    .y(log_smally),
    .cin(nsrcin),
    .r(log_small_adder_n733));
  /* fppow16.vhdl:3340:35  */
  assign n737 = log_small[22]; // extract
  /* fppow16.vhdl:3340:21  */
  assign n738 = n737 ? 2'b11 : n743;
  /* fppow16.vhdl:3341:35  */
  assign n740 = log_small[22:21]; // extract
  /* fppow16.vhdl:3341:56  */
  assign n742 = n740 == 2'b01;
  /* fppow16.vhdl:3341:11  */
  assign n743 = n742 ? 2'b10 : 2'b01;
  /* fppow16.vhdl:3346:47  */
  assign n746 = {4'b0011, e0_sub};
  /* fppow16.vhdl:3346:66  */
  assign n748 = {1'b0, lzo_d3};
  /* fppow16.vhdl:3346:58  */
  assign n749 = n746 - n748;
  /* fppow16.vhdl:3347:18  */
  assign n750 = e_small[5]; // extract
  /* fppow16.vhdl:3348:32  */
  assign n751 = log_small[22:2]; // extract
  /* fppow16.vhdl:3348:64  */
  assign n752 = log_small[22]; // extract
  /* fppow16.vhdl:3348:50  */
  assign n753 = n752 ? n751 : n756;
  /* fppow16.vhdl:3349:26  */
  assign n754 = log_small[21:1]; // extract
  /* fppow16.vhdl:3349:57  */
  assign n755 = log_small[21]; // extract
  /* fppow16.vhdl:3349:12  */
  assign n756 = n755 ? n754 : n757;
  /* fppow16.vhdl:3350:26  */
  assign n757 = log_small[20:0]; // extract
  /* fppow16.vhdl:3352:20  */
  assign n759 = e_small_d3[4:0]; // extract
  /* fppow16.vhdl:3352:33  */
  assign n760 = small_d5 ? n759 : n763;
  /* fppow16.vhdl:3353:47  */
  assign n762 = {1'b0, e_normal};
  /* fppow16.vhdl:3353:24  */
  assign n763 = e0offset_d9 - n762;
  /* fppow16.vhdl:3354:32  */
  assign n764 = log_small_normd_d3[19:0]; // extract
  /* fppow16.vhdl:3354:50  */
  assign n766 = {n764, 1'b0};
  /* fppow16.vhdl:3354:56  */
  assign n767 = small_d5 ? n766 : n768;
  /* fppow16.vhdl:3355:28  */
  assign n768 = log_normal_normd[28:8]; // extract
  /* fppow16.vhdl:3356:18  */
  assign n769 = log_g[3]; // extract
  /* fppow16.vhdl:3358:23  */
  assign n770 = log_g[20:4]; // extract
  /* fppow16.vhdl:3358:16  */
  assign n771 = {er, n770};
  /* fppow16.vhdl:3359:39  */
  assign n773 = {21'b000000000000000000000, round};
  /* fppow16.vhdl:3360:4  */
  intadder_22_freq500_uid55 finalroundadder (
    .clk(clk),
    .x(frax),
    .y(fray),
    .cin(n774),
    .r(finalroundadder_n775));
  /* fppow16.vhdl:3366:36  */
  assign n779 = xexnsgn_d10[2]; // extract
  /* fppow16.vhdl:3366:56  */
  assign n780 = xexnsgn_d10[1]; // extract
  /* fppow16.vhdl:3366:74  */
  assign n781 = xexnsgn_d10[0]; // extract
  /* fppow16.vhdl:3366:60  */
  assign n782 = n780 | n781;
  /* fppow16.vhdl:3366:40  */
  assign n783 = n779 & n782;
  /* fppow16.vhdl:3366:95  */
  assign n784 = xexnsgn_d10[1]; // extract
  /* fppow16.vhdl:3366:114  */
  assign n785 = xexnsgn_d10[0]; // extract
  /* fppow16.vhdl:3366:99  */
  assign n786 = n784 & n785;
  /* fppow16.vhdl:3366:80  */
  assign n787 = n783 | n786;
  /* fppow16.vhdl:3366:18  */
  assign n788 = n787 ? 3'b110 : n793;
  /* fppow16.vhdl:3367:53  */
  assign n790 = xexnsgn_d10[2:1]; // extract
  /* fppow16.vhdl:3367:66  */
  assign n792 = n790 == 2'b00;
  /* fppow16.vhdl:3366:126  */
  assign n793 = n792 ? 3'b101 : n798;
  /* fppow16.vhdl:3368:53  */
  assign n795 = xexnsgn_d10[2:1]; // extract
  /* fppow16.vhdl:3368:66  */
  assign n797 = n795 == 2'b10;
  /* fppow16.vhdl:3367:74  */
  assign n798 = n797 ? 3'b100 : n811;
  /* fppow16.vhdl:3369:36  */
  assign n800 = {2'b00, sr_d10};
  /* fppow16.vhdl:3369:72  */
  assign n801 = log_normal_normd_d1[29]; // extract
  /* fppow16.vhdl:3369:86  */
  assign n802 = ~n801;
  /* fppow16.vhdl:3369:105  */
  assign n803 = ~small_d6;
  /* fppow16.vhdl:3369:92  */
  assign n804 = n803 & n802;
  /* fppow16.vhdl:3369:137  */
  assign n805 = log_small_normd_d4[20]; // extract
  /* fppow16.vhdl:3369:145  */
  assign n806 = ~n805;
  /* fppow16.vhdl:3369:151  */
  assign n807 = small_d6 & n806;
  /* fppow16.vhdl:3369:112  */
  assign n808 = n804 | n807;
  /* fppow16.vhdl:3369:189  */
  assign n809 = small_d6 & ufl_d4;
  /* fppow16.vhdl:3369:172  */
  assign n810 = n808 | n809;
  /* fppow16.vhdl:3368:74  */
  assign n811 = n810 ? n800 : n813;
  /* fppow16.vhdl:3370:37  */
  assign n813 = {2'b01, sr_d10};
  /* fppow16.vhdl:3371:14  */
  assign n814 = {rexn, efr};
  /* fppow16.vhdl:3132:10  */
  always @(posedge clk)
    n815 <= xexnsgn;
  /* fppow16.vhdl:3132:10  */
  always @(posedge clk)
    n816 <= xexnsgn_d1;
  /* fppow16.vhdl:3132:10  */
  always @(posedge clk)
    n817 <= xexnsgn_d2;
  /* fppow16.vhdl:3132:10  */
  always @(posedge clk)
    n818 <= xexnsgn_d3;
  /* fppow16.vhdl:3132:10  */
  always @(posedge clk)
    n819 <= xexnsgn_d4;
  /* fppow16.vhdl:3132:10  */
  always @(posedge clk)
    n820 <= xexnsgn_d5;
  /* fppow16.vhdl:3132:10  */
  always @(posedge clk)
    n821 <= xexnsgn_d6;
  /* fppow16.vhdl:3132:10  */
  always @(posedge clk)
    n822 <= xexnsgn_d7;
  /* fppow16.vhdl:3132:10  */
  always @(posedge clk)
    n823 <= xexnsgn_d8;
  /* fppow16.vhdl:3132:10  */
  always @(posedge clk)
    n824 <= xexnsgn_d9;
  /* fppow16.vhdl:3132:10  */
  always @(posedge clk)
    n825 <= y0;
  /* fppow16.vhdl:3132:10  */
  always @(posedge clk)
    n826 <= sr;
  /* fppow16.vhdl:3132:10  */
  always @(posedge clk)
    n827 <= sr_d1;
  /* fppow16.vhdl:3132:10  */
  always @(posedge clk)
    n828 <= sr_d2;
  /* fppow16.vhdl:3132:10  */
  always @(posedge clk)
    n829 <= sr_d3;
  /* fppow16.vhdl:3132:10  */
  always @(posedge clk)
    n830 <= sr_d4;
  /* fppow16.vhdl:3132:10  */
  always @(posedge clk)
    n831 <= sr_d5;
  /* fppow16.vhdl:3132:10  */
  always @(posedge clk)
    n832 <= sr_d6;
  /* fppow16.vhdl:3132:10  */
  always @(posedge clk)
    n833 <= sr_d7;
  /* fppow16.vhdl:3132:10  */
  always @(posedge clk)
    n834 <= sr_d8;
  /* fppow16.vhdl:3132:10  */
  always @(posedge clk)
    n835 <= sr_d9;
  /* fppow16.vhdl:3132:10  */
  always @(posedge clk)
    n836 <= eeqzero;
  /* fppow16.vhdl:3132:10  */
  always @(posedge clk)
    n837 <= eeqzero_d1;
  /* fppow16.vhdl:3132:10  */
  always @(posedge clk)
    n838 <= eeqzero_d2;
  /* fppow16.vhdl:3132:10  */
  always @(posedge clk)
    n839 <= eeqzero_d3;
  /* fppow16.vhdl:3132:10  */
  always @(posedge clk)
    n840 <= lzo;
  /* fppow16.vhdl:3132:10  */
  always @(posedge clk)
    n841 <= lzo_d1;
  /* fppow16.vhdl:3132:10  */
  always @(posedge clk)
    n842 <= lzo_d2;
  /* fppow16.vhdl:3132:10  */
  always @(posedge clk)
    n843 <= pfinal_s;
  /* fppow16.vhdl:3132:10  */
  always @(posedge clk)
    n844 <= pfinal_s_d1;
  /* fppow16.vhdl:3132:10  */
  always @(posedge clk)
    n845 <= pfinal_s_d2;
  /* fppow16.vhdl:3132:10  */
  always @(posedge clk)
    n846 <= dorr;
  /* fppow16.vhdl:3132:10  */
  always @(posedge clk)
    n847 <= dorr_d1;
  /* fppow16.vhdl:3132:10  */
  always @(posedge clk)
    n848 <= \small ;
  /* fppow16.vhdl:3132:10  */
  always @(posedge clk)
    n849 <= small_d1;
  /* fppow16.vhdl:3132:10  */
  always @(posedge clk)
    n850 <= small_d2;
  /* fppow16.vhdl:3132:10  */
  always @(posedge clk)
    n851 <= small_d3;
  /* fppow16.vhdl:3132:10  */
  always @(posedge clk)
    n852 <= small_d4;
  /* fppow16.vhdl:3132:10  */
  always @(posedge clk)
    n853 <= small_d5;
  /* fppow16.vhdl:3132:10  */
  always @(posedge clk)
    n854 <= small_absz0_normd;
  /* fppow16.vhdl:3132:10  */
  always @(posedge clk)
    n855 <= inva0;
  /* fppow16.vhdl:3132:10  */
  always @(posedge clk)
    n856 <= a1;
  /* fppow16.vhdl:3132:10  */
  always @(posedge clk)
    n857 <= zm1;
  /* fppow16.vhdl:3132:10  */
  always @(posedge clk)
    n858 <= zfinal;
  /* fppow16.vhdl:3132:10  */
  always @(posedge clk)
    n859 <= zfinal_d1;
  /* fppow16.vhdl:3132:10  */
  always @(posedge clk)
    n860 <= log_normal_normd;
  /* fppow16.vhdl:3132:10  */
  always @(posedge clk)
    n861 <= e_small;
  /* fppow16.vhdl:3132:10  */
  always @(posedge clk)
    n862 <= e_small_d1;
  /* fppow16.vhdl:3132:10  */
  always @(posedge clk)
    n863 <= e_small_d2;
  /* fppow16.vhdl:3132:10  */
  always @(posedge clk)
    n864 <= ufl;
  /* fppow16.vhdl:3132:10  */
  always @(posedge clk)
    n865 <= ufl_d1;
  /* fppow16.vhdl:3132:10  */
  always @(posedge clk)
    n866 <= ufl_d2;
  /* fppow16.vhdl:3132:10  */
  always @(posedge clk)
    n867 <= ufl_d3;
  /* fppow16.vhdl:3132:10  */
  always @(posedge clk)
    n868 <= log_small_normd;
  /* fppow16.vhdl:3132:10  */
  always @(posedge clk)
    n869 <= log_small_normd_d1;
  /* fppow16.vhdl:3132:10  */
  always @(posedge clk)
    n870 <= log_small_normd_d2;
  /* fppow16.vhdl:3132:10  */
  always @(posedge clk)
    n871 <= log_small_normd_d3;
  /* fppow16.vhdl:3132:10  */
  always @(posedge clk)
    n872 <= e0offset;
  /* fppow16.vhdl:3132:10  */
  always @(posedge clk)
    n873 <= e0offset_d1;
  /* fppow16.vhdl:3132:10  */
  always @(posedge clk)
    n874 <= e0offset_d2;
  /* fppow16.vhdl:3132:10  */
  always @(posedge clk)
    n875 <= e0offset_d3;
  /* fppow16.vhdl:3132:10  */
  always @(posedge clk)
    n876 <= e0offset_d4;
  /* fppow16.vhdl:3132:10  */
  always @(posedge clk)
    n877 <= e0offset_d5;
  /* fppow16.vhdl:3132:10  */
  always @(posedge clk)
    n878 <= e0offset_d6;
  /* fppow16.vhdl:3132:10  */
  always @(posedge clk)
    n879 <= e0offset_d7;
  /* fppow16.vhdl:3132:10  */
  always @(posedge clk)
    n880 <= e0offset_d8;
endmodule

module lzc_10_freq500_uid7
  (input  clk,
   input  [9:0] i,
   output [3:0] o);
  wire [14:0] level4;
  wire digit3;
  wire [6:0] level3;
  wire [6:0] level3_d1;
  wire digit2;
  wire digit2_d1;
  wire [2:0] level2;
  wire [1:0] lowbits;
  wire [1:0] outhighbits;
  wire [1:0] outhighbits_d1;
  wire [14:0] n458;
  wire [7:0] n460;
  wire n462;
  wire n463;
  wire [6:0] n465;
  wire [6:0] n466;
  wire [6:0] n467;
  wire [3:0] n469;
  wire n471;
  wire n472;
  wire [2:0] n474;
  wire [2:0] n475;
  wire [2:0] n476;
  wire n479;
  wire n482;
  wire n485;
  wire n488;
  wire [3:0] n490;
  reg [1:0] n491;
  wire [1:0] n492;
  wire [3:0] n494;
  reg [6:0] n495;
  reg n496;
  reg [1:0] n497;
  assign o = n494; //(module output)
  /* fppow16.vhdl:1854:8  */
  assign level4 = n458; // (signal)
  /* fppow16.vhdl:1856:8  */
  assign digit3 = n463; // (signal)
  /* fppow16.vhdl:1858:8  */
  assign level3 = n466; // (signal)
  /* fppow16.vhdl:1858:16  */
  assign level3_d1 = n495; // (signal)
  /* fppow16.vhdl:1860:8  */
  assign digit2 = n472; // (signal)
  /* fppow16.vhdl:1860:16  */
  assign digit2_d1 = n496; // (signal)
  /* fppow16.vhdl:1862:8  */
  assign level2 = n475; // (signal)
  /* fppow16.vhdl:1864:8  */
  assign lowbits = n491; // (signal)
  /* fppow16.vhdl:1866:8  */
  assign outhighbits = n492; // (signal)
  /* fppow16.vhdl:1866:21  */
  assign outhighbits_d1 = n497; // (signal)
  /* fppow16.vhdl:1878:16  */
  assign n458 = {i, 5'b11111};
  /* fppow16.vhdl:1880:28  */
  assign n460 = level4[14:7]; // extract
  /* fppow16.vhdl:1880:42  */
  assign n462 = n460 == 8'b00000000;
  /* fppow16.vhdl:1880:17  */
  assign n463 = n462 ? 1'b1 : 1'b0;
  /* fppow16.vhdl:1881:19  */
  assign n465 = level4[6:0]; // extract
  /* fppow16.vhdl:1881:32  */
  assign n466 = digit3 ? n465 : n467;
  /* fppow16.vhdl:1881:59  */
  assign n467 = level4[14:8]; // extract
  /* fppow16.vhdl:1882:28  */
  assign n469 = level3[6:3]; // extract
  /* fppow16.vhdl:1882:41  */
  assign n471 = n469 == 4'b0000;
  /* fppow16.vhdl:1882:17  */
  assign n472 = n471 ? 1'b1 : 1'b0;
  /* fppow16.vhdl:1883:22  */
  assign n474 = level3_d1[2:0]; // extract
  /* fppow16.vhdl:1883:35  */
  assign n475 = digit2_d1 ? n474 : n476;
  /* fppow16.vhdl:1883:68  */
  assign n476 = level3_d1[6:4]; // extract
  /* fppow16.vhdl:1886:12  */
  assign n479 = level2 == 3'b000;
  /* fppow16.vhdl:1887:12  */
  assign n482 = level2 == 3'b001;
  /* fppow16.vhdl:1888:12  */
  assign n485 = level2 == 3'b010;
  /* fppow16.vhdl:1889:12  */
  assign n488 = level2 == 3'b011;
  assign n490 = {n488, n485, n482, n479};
  /* fppow16.vhdl:1885:4  */
  always @*
    case (n490)
      4'b1000: n491 = 2'b01;
      4'b0100: n491 = 2'b01;
      4'b0010: n491 = 2'b10;
      4'b0001: n491 = 2'b11;
      default: n491 = 2'b00;
    endcase
  /* fppow16.vhdl:1891:35  */
  assign n492 = {digit3, digit2};
  /* fppow16.vhdl:1892:24  */
  assign n494 = {outhighbits_d1, lowbits};
  /* fppow16.vhdl:1871:10  */
  always @(posedge clk)
    n495 <= level3;
  /* fppow16.vhdl:1871:10  */
  always @(posedge clk)
    n496 <= digit2;
  /* fppow16.vhdl:1871:10  */
  always @(posedge clk)
    n497 <= outhighbits;
endmodule

module intadder_16_freq500_uid5
  (input  clk,
   input  [15:0] x,
   input  [15:0] y,
   input  cin,
   output [15:0] r);
  wire [15:0] rtmp;
  wire [15:0] n446;
  wire [15:0] n447;
  wire [15:0] n448;
  assign r = rtmp; //(module output)
  /* fppow16.vhdl:1817:8  */
  assign rtmp = n448; // (signal)
  /* fppow16.vhdl:1820:14  */
  assign n446 = x + y;
  /* fppow16.vhdl:1820:18  */
  assign n447 = {15'b0, cin};  //  uext
  /* fppow16.vhdl:1820:18  */
  assign n448 = n446 + n447;
endmodule

module top_module
  (input  clk,
   input  [17:0] X,
   input  [17:0] Y,
   output [17:0] R);
  wire [1:0] flagsx;
  wire signx;
  wire signx_d1;
  wire signx_d2;
  wire [4:0] expfieldx;
  wire [9:0] fracx;
  wire [1:0] flagsy;
  wire signy;
  wire signy_d1;
  wire signy_d2;
  wire signy_d3;
  wire [4:0] expfieldy;
  wire [9:0] fracy;
  wire zerox;
  wire zerox_d1;
  wire zerox_d2;
  wire zerox_d3;
  wire zeroy;
  wire zeroy_d1;
  wire zeroy_d2;
  wire normalx;
  wire normalx_d1;
  wire normalx_d2;
  wire normaly;
  wire normaly_d1;
  wire normaly_d2;
  wire normaly_d3;
  wire infx;
  wire infx_d1;
  wire infx_d2;
  wire infx_d3;
  wire infy;
  wire infy_d1;
  wire infy_d2;
  wire infy_d3;
  wire s_nan_in;
  wire s_nan_in_d1;
  wire s_nan_in_d2;
  wire [14:0] oneexpfrac;
  wire [15:0] expfracx;
  wire [15:0] oneexpfraccompl;
  wire [15:0] cmpxoneres;
  wire xisoneandnormal;
  wire absxgtoneandnormal;
  wire absxgtoneandnormal_d1;
  wire absxgtoneandnormal_d2;
  wire absxgtoneandnormal_d3;
  wire absxltoneandnormal;
  wire absxltoneandnormal_d1;
  wire absxltoneandnormal_d2;
  wire absxltoneandnormal_d3;
  wire [9:0] fracyreverted;
  wire [3:0] z_righty;
  wire [3:0] z_righty_d1;
  wire [5:0] weightlsbypre;
  wire [5:0] weightlsbypre_d1;
  wire [5:0] weightlsbypre_d2;
  wire [5:0] weightlsby;
  wire oddinty;
  wire oddinty_d1;
  wire eveninty;
  wire eveninty_d1;
  wire notintnormaly;
  wire risinfspecialcase;
  wire risinfspecialcase_d1;
  wire risinfspecialcase_d2;
  wire risinfspecialcase_d3;
  wire risinfspecialcase_d4;
  wire risinfspecialcase_d5;
  wire risinfspecialcase_d6;
  wire risinfspecialcase_d7;
  wire risinfspecialcase_d8;
  wire risinfspecialcase_d9;
  wire risinfspecialcase_d10;
  wire risinfspecialcase_d11;
  wire risinfspecialcase_d12;
  wire risinfspecialcase_d13;
  wire risinfspecialcase_d14;
  wire risinfspecialcase_d15;
  wire risinfspecialcase_d16;
  wire riszerospecialcase;
  wire riszerospecialcase_d1;
  wire riszerospecialcase_d2;
  wire riszerospecialcase_d3;
  wire riszerospecialcase_d4;
  wire riszerospecialcase_d5;
  wire riszerospecialcase_d6;
  wire riszerospecialcase_d7;
  wire riszerospecialcase_d8;
  wire riszerospecialcase_d9;
  wire riszerospecialcase_d10;
  wire riszerospecialcase_d11;
  wire riszerospecialcase_d12;
  wire riszerospecialcase_d13;
  wire riszerospecialcase_d14;
  wire riszerospecialcase_d15;
  wire riszerospecialcase_d16;
  wire risone;
  wire risone_d1;
  wire risone_d2;
  wire risone_d3;
  wire risone_d4;
  wire risone_d5;
  wire risone_d6;
  wire risone_d7;
  wire risone_d8;
  wire risone_d9;
  wire risone_d10;
  wire risone_d11;
  wire risone_d12;
  wire risone_d13;
  wire risone_d14;
  wire risone_d15;
  wire risone_d16;
  wire risone_d17;
  wire risone_d18;
  wire risone_d19;
  wire risnan;
  wire risnan_d1;
  wire risnan_d2;
  wire risnan_d3;
  wire risnan_d4;
  wire risnan_d5;
  wire risnan_d6;
  wire risnan_d7;
  wire risnan_d8;
  wire risnan_d9;
  wire risnan_d10;
  wire risnan_d11;
  wire risnan_d12;
  wire risnan_d13;
  wire risnan_d14;
  wire risnan_d15;
  wire risnan_d16;
  wire risnan_d17;
  wire signr;
  wire signr_d1;
  wire signr_d2;
  wire signr_d3;
  wire signr_d4;
  wire signr_d5;
  wire signr_d6;
  wire signr_d7;
  wire signr_d8;
  wire signr_d9;
  wire signr_d10;
  wire signr_d11;
  wire signr_d12;
  wire signr_d13;
  wire signr_d14;
  wire signr_d15;
  wire signr_d16;
  wire signr_d17;
  wire [24:0] login;
  wire [24:0] lnx;
  wire [25:0] p;
  wire [17:0] e;
  wire [17:0] e_d1;
  wire [1:0] flagse;
  wire [1:0] flagse_d1;
  wire riszerofromexp;
  wire riszero;
  wire risinffromexp;
  wire risinf;
  wire [1:0] flagr;
  wire [14:0] r_expfrac;
  wire [1:0] n126;
  wire n127;
  wire [4:0] n128;
  wire [9:0] n129;
  wire [1:0] n130;
  wire n131;
  wire [4:0] n132;
  wire [9:0] n133;
  wire n136;
  wire n137;
  wire n141;
  wire n142;
  wire n146;
  wire n147;
  wire n151;
  wire n152;
  wire n156;
  wire n157;
  wire n161;
  wire n162;
  wire n166;
  wire n168;
  wire n169;
  wire n170;
  wire [5:0] n174;
  wire [15:0] n175;
  wire [14:0] n176;
  wire [15:0] n178;
  localparam n179 = 1'b1;
  wire [15:0] cmpxone_n180;
  wire [17:0] n185;
  wire n186;
  wire n187;
  wire n189;
  wire n190;
  wire n191;
  wire n192;
  wire n193;
  wire n194;
  wire n195;
  wire n196;
  wire n197;
  wire [1:0] n198;
  wire n199;
  wire [2:0] n200;
  wire n201;
  wire [3:0] n202;
  wire n203;
  wire [4:0] n204;
  wire n205;
  wire [5:0] n206;
  wire n207;
  wire [6:0] n208;
  wire n209;
  wire [7:0] n210;
  wire n211;
  wire [8:0] n212;
  wire n213;
  wire [9:0] n214;
  wire [3:0] fppow_5_10_freq500_uid2right1counter_n215;
  wire [5:0] n219;
  wire [5:0] n221;
  wire [5:0] n222;
  wire [5:0] n223;
  wire n225;
  wire n226;
  wire n228;
  wire n229;
  wire n230;
  wire n231;
  wire n232;
  wire n234;
  wire n235;
  wire n237;
  wire n238;
  wire n239;
  wire n240;
  wire n241;
  wire n242;
  wire n243;
  wire n244;
  wire n245;
  wire n246;
  wire n247;
  wire n248;
  wire n249;
  wire n250;
  wire n251;
  wire n252;
  wire n253;
  wire n254;
  wire n255;
  wire n256;
  wire n257;
  wire n258;
  wire n259;
  wire n260;
  wire n261;
  wire n262;
  wire n263;
  wire n264;
  wire n265;
  wire n266;
  wire n267;
  wire n268;
  wire n269;
  wire n270;
  wire n271;
  wire n272;
  wire n273;
  wire n274;
  wire n275;
  wire n276;
  wire n277;
  wire n278;
  wire n279;
  wire n280;
  wire n281;
  wire n282;
  wire n283;
  wire [2:0] n285;
  wire [7:0] n286;
  wire [17:0] n287;
  wire [24:0] n289;
  wire [24:0] fppow_5_10_freq500_uid2log_n290;
  wire [25:0] fppow_5_10_freq500_uid2mult_n293;
  wire [17:0] fppow_5_10_freq500_uid2exp_n296;
  wire [1:0] n299;
  wire n302;
  wire n303;
  wire n305;
  wire n308;
  wire n309;
  wire n311;
  wire [1:0] n313;
  wire [1:0] n315;
  wire [1:0] n317;
  wire [14:0] n320;
  wire [14:0] n321;
  wire [2:0] n322;
  wire [17:0] n323;
  reg n324;
  reg n325;
  reg n326;
  reg n327;
  reg n328;
  reg n329;
  reg n330;
  reg n331;
  reg n332;
  reg n333;
  reg n334;
  reg n335;
  reg n336;
  reg n337;
  reg n338;
  reg n339;
  reg n340;
  reg n341;
  reg n342;
  reg n343;
  reg n344;
  reg n345;
  reg n346;
  reg n347;
  reg n348;
  reg n349;
  reg n350;
  reg n351;
  reg n352;
  reg [3:0] n353;
  reg [5:0] n354;
  reg [5:0] n355;
  reg n356;
  reg n357;
  reg n358;
  reg n359;
  reg n360;
  reg n361;
  reg n362;
  reg n363;
  reg n364;
  reg n365;
  reg n366;
  reg n367;
  reg n368;
  reg n369;
  reg n370;
  reg n371;
  reg n372;
  reg n373;
  reg n374;
  reg n375;
  reg n376;
  reg n377;
  reg n378;
  reg n379;
  reg n380;
  reg n381;
  reg n382;
  reg n383;
  reg n384;
  reg n385;
  reg n386;
  reg n387;
  reg n388;
  reg n389;
  reg n390;
  reg n391;
  reg n392;
  reg n393;
  reg n394;
  reg n395;
  reg n396;
  reg n397;
  reg n398;
  reg n399;
  reg n400;
  reg n401;
  reg n402;
  reg n403;
  reg n404;
  reg n405;
  reg n406;
  reg n407;
  reg n408;
  reg n409;
  reg n410;
  reg n411;
  reg n412;
  reg n413;
  reg n414;
  reg n415;
  reg n416;
  reg n417;
  reg n418;
  reg n419;
  reg n420;
  reg n421;
  reg n422;
  reg n423;
  reg n424;
  reg n425;
  reg n426;
  reg n427;
  reg n428;
  reg n429;
  reg n430;
  reg n431;
  reg n432;
  reg n433;
  reg n434;
  reg n435;
  reg n436;
  reg n437;
  reg n438;
  reg n439;
  reg n440;
  reg n441;
  reg n442;
  reg [17:0] n443;
  reg [1:0] n444;
  assign R = n323; //(module output)
  /* fppow16.vhdl:4920:8  */
  assign flagsx = n126; // (signal)
  /* fppow16.vhdl:4922:8  */
  assign signx = n127; // (signal)
  /* fppow16.vhdl:4922:15  */
  assign signx_d1 = n324; // (signal)
  /* fppow16.vhdl:4922:25  */
  assign signx_d2 = n325; // (signal)
  /* fppow16.vhdl:4924:8  */
  assign expfieldx = n128; // (signal)
  /* fppow16.vhdl:4926:8  */
  assign fracx = n129; // (signal)
  /* fppow16.vhdl:4928:8  */
  assign flagsy = n130; // (signal)
  /* fppow16.vhdl:4930:8  */
  assign signy = n131; // (signal)
  /* fppow16.vhdl:4930:15  */
  assign signy_d1 = n326; // (signal)
  /* fppow16.vhdl:4930:25  */
  assign signy_d2 = n327; // (signal)
  /* fppow16.vhdl:4930:35  */
  assign signy_d3 = n328; // (signal)
  /* fppow16.vhdl:4932:8  */
  assign expfieldy = n132; // (signal)
  /* fppow16.vhdl:4934:8  */
  assign fracy = n133; // (signal)
  /* fppow16.vhdl:4936:8  */
  assign zerox = n137; // (signal)
  /* fppow16.vhdl:4936:15  */
  assign zerox_d1 = n329; // (signal)
  /* fppow16.vhdl:4936:25  */
  assign zerox_d2 = n330; // (signal)
  /* fppow16.vhdl:4936:35  */
  assign zerox_d3 = n331; // (signal)
  /* fppow16.vhdl:4938:8  */
  assign zeroy = n142; // (signal)
  /* fppow16.vhdl:4938:15  */
  assign zeroy_d1 = n332; // (signal)
  /* fppow16.vhdl:4938:25  */
  assign zeroy_d2 = n333; // (signal)
  /* fppow16.vhdl:4940:8  */
  assign normalx = n147; // (signal)
  /* fppow16.vhdl:4940:17  */
  assign normalx_d1 = n334; // (signal)
  /* fppow16.vhdl:4940:29  */
  assign normalx_d2 = n335; // (signal)
  /* fppow16.vhdl:4942:8  */
  assign normaly = n152; // (signal)
  /* fppow16.vhdl:4942:17  */
  assign normaly_d1 = n336; // (signal)
  /* fppow16.vhdl:4942:29  */
  assign normaly_d2 = n337; // (signal)
  /* fppow16.vhdl:4942:41  */
  assign normaly_d3 = n338; // (signal)
  /* fppow16.vhdl:4944:8  */
  assign infx = n157; // (signal)
  /* fppow16.vhdl:4944:14  */
  assign infx_d1 = n339; // (signal)
  /* fppow16.vhdl:4944:23  */
  assign infx_d2 = n340; // (signal)
  /* fppow16.vhdl:4944:32  */
  assign infx_d3 = n341; // (signal)
  /* fppow16.vhdl:4946:8  */
  assign infy = n162; // (signal)
  /* fppow16.vhdl:4946:14  */
  assign infy_d1 = n342; // (signal)
  /* fppow16.vhdl:4946:23  */
  assign infy_d2 = n343; // (signal)
  /* fppow16.vhdl:4946:32  */
  assign infy_d3 = n344; // (signal)
  /* fppow16.vhdl:4948:8  */
  assign s_nan_in = n170; // (signal)
  /* fppow16.vhdl:4948:18  */
  assign s_nan_in_d1 = n345; // (signal)
  /* fppow16.vhdl:4948:31  */
  assign s_nan_in_d2 = n346; // (signal)
  /* fppow16.vhdl:4950:8  */
  assign oneexpfrac = 15'b011110000000000; // (signal)
  /* fppow16.vhdl:4952:8  */
  assign expfracx = n175; // (signal)
  /* fppow16.vhdl:4954:8  */
  assign oneexpfraccompl = n178; // (signal)
  /* fppow16.vhdl:4956:8  */
  assign cmpxoneres = cmpxone_n180; // (signal)
  /* fppow16.vhdl:4958:8  */
  assign xisoneandnormal = n187; // (signal)
  /* fppow16.vhdl:4960:8  */
  assign absxgtoneandnormal = n193; // (signal)
  /* fppow16.vhdl:4960:28  */
  assign absxgtoneandnormal_d1 = n347; // (signal)
  /* fppow16.vhdl:4960:51  */
  assign absxgtoneandnormal_d2 = n348; // (signal)
  /* fppow16.vhdl:4960:74  */
  assign absxgtoneandnormal_d3 = n349; // (signal)
  /* fppow16.vhdl:4962:8  */
  assign absxltoneandnormal = n195; // (signal)
  /* fppow16.vhdl:4962:28  */
  assign absxltoneandnormal_d1 = n350; // (signal)
  /* fppow16.vhdl:4962:51  */
  assign absxltoneandnormal_d2 = n351; // (signal)
  /* fppow16.vhdl:4962:74  */
  assign absxltoneandnormal_d3 = n352; // (signal)
  /* fppow16.vhdl:4964:8  */
  assign fracyreverted = n214; // (signal)
  /* fppow16.vhdl:4966:8  */
  assign z_righty = fppow_5_10_freq500_uid2right1counter_n215; // (signal)
  /* fppow16.vhdl:4966:18  */
  assign z_righty_d1 = n353; // (signal)
  /* fppow16.vhdl:4968:8  */
  assign weightlsbypre = n221; // (signal)
  /* fppow16.vhdl:4968:23  */
  assign weightlsbypre_d1 = n354; // (signal)
  /* fppow16.vhdl:4968:41  */
  assign weightlsbypre_d2 = n355; // (signal)
  /* fppow16.vhdl:4970:8  */
  assign weightlsby = n223; // (signal)
  /* fppow16.vhdl:4972:8  */
  assign oddinty = n226; // (signal)
  /* fppow16.vhdl:4972:17  */
  assign oddinty_d1 = n356; // (signal)
  /* fppow16.vhdl:4974:8  */
  assign eveninty = n232; // (signal)
  /* fppow16.vhdl:4974:18  */
  assign eveninty_d1 = n357; // (signal)
  /* fppow16.vhdl:4976:8  */
  assign notintnormaly = n235; // (signal)
  /* fppow16.vhdl:4978:8  */
  assign risinfspecialcase = n253; // (signal)
  /* fppow16.vhdl:4978:27  */
  assign risinfspecialcase_d1 = n358; // (signal)
  /* fppow16.vhdl:4978:49  */
  assign risinfspecialcase_d2 = n359; // (signal)
  /* fppow16.vhdl:4978:71  */
  assign risinfspecialcase_d3 = n360; // (signal)
  /* fppow16.vhdl:4978:93  */
  assign risinfspecialcase_d4 = n361; // (signal)
  /* fppow16.vhdl:4978:115  */
  assign risinfspecialcase_d5 = n362; // (signal)
  /* fppow16.vhdl:4978:137  */
  assign risinfspecialcase_d6 = n363; // (signal)
  /* fppow16.vhdl:4978:159  */
  assign risinfspecialcase_d7 = n364; // (signal)
  /* fppow16.vhdl:4978:181  */
  assign risinfspecialcase_d8 = n365; // (signal)
  /* fppow16.vhdl:4978:203  */
  assign risinfspecialcase_d9 = n366; // (signal)
  /* fppow16.vhdl:4978:225  */
  assign risinfspecialcase_d10 = n367; // (signal)
  /* fppow16.vhdl:4978:248  */
  assign risinfspecialcase_d11 = n368; // (signal)
  /* fppow16.vhdl:4978:271  */
  assign risinfspecialcase_d12 = n369; // (signal)
  /* fppow16.vhdl:4978:294  */
  assign risinfspecialcase_d13 = n370; // (signal)
  /* fppow16.vhdl:4978:317  */
  assign risinfspecialcase_d14 = n371; // (signal)
  /* fppow16.vhdl:4978:340  */
  assign risinfspecialcase_d15 = n372; // (signal)
  /* fppow16.vhdl:4978:363  */
  assign risinfspecialcase_d16 = n373; // (signal)
  /* fppow16.vhdl:4980:8  */
  assign riszerospecialcase = n271; // (signal)
  /* fppow16.vhdl:4980:28  */
  assign riszerospecialcase_d1 = n374; // (signal)
  /* fppow16.vhdl:4980:51  */
  assign riszerospecialcase_d2 = n375; // (signal)
  /* fppow16.vhdl:4980:74  */
  assign riszerospecialcase_d3 = n376; // (signal)
  /* fppow16.vhdl:4980:97  */
  assign riszerospecialcase_d4 = n377; // (signal)
  /* fppow16.vhdl:4980:120  */
  assign riszerospecialcase_d5 = n378; // (signal)
  /* fppow16.vhdl:4980:143  */
  assign riszerospecialcase_d6 = n379; // (signal)
  /* fppow16.vhdl:4980:166  */
  assign riszerospecialcase_d7 = n380; // (signal)
  /* fppow16.vhdl:4980:189  */
  assign riszerospecialcase_d8 = n381; // (signal)
  /* fppow16.vhdl:4980:212  */
  assign riszerospecialcase_d9 = n382; // (signal)
  /* fppow16.vhdl:4980:235  */
  assign riszerospecialcase_d10 = n383; // (signal)
  /* fppow16.vhdl:4980:259  */
  assign riszerospecialcase_d11 = n384; // (signal)
  /* fppow16.vhdl:4980:283  */
  assign riszerospecialcase_d12 = n385; // (signal)
  /* fppow16.vhdl:4980:307  */
  assign riszerospecialcase_d13 = n386; // (signal)
  /* fppow16.vhdl:4980:331  */
  assign riszerospecialcase_d14 = n387; // (signal)
  /* fppow16.vhdl:4980:355  */
  assign riszerospecialcase_d15 = n388; // (signal)
  /* fppow16.vhdl:4980:379  */
  assign riszerospecialcase_d16 = n389; // (signal)
  /* fppow16.vhdl:4982:8  */
  assign risone = n277; // (signal)
  /* fppow16.vhdl:4982:16  */
  assign risone_d1 = n390; // (signal)
  /* fppow16.vhdl:4982:27  */
  assign risone_d2 = n391; // (signal)
  /* fppow16.vhdl:4982:38  */
  assign risone_d3 = n392; // (signal)
  /* fppow16.vhdl:4982:49  */
  assign risone_d4 = n393; // (signal)
  /* fppow16.vhdl:4982:60  */
  assign risone_d5 = n394; // (signal)
  /* fppow16.vhdl:4982:71  */
  assign risone_d6 = n395; // (signal)
  /* fppow16.vhdl:4982:82  */
  assign risone_d7 = n396; // (signal)
  /* fppow16.vhdl:4982:93  */
  assign risone_d8 = n397; // (signal)
  /* fppow16.vhdl:4982:104  */
  assign risone_d9 = n398; // (signal)
  /* fppow16.vhdl:4982:115  */
  assign risone_d10 = n399; // (signal)
  /* fppow16.vhdl:4982:127  */
  assign risone_d11 = n400; // (signal)
  /* fppow16.vhdl:4982:139  */
  assign risone_d12 = n401; // (signal)
  /* fppow16.vhdl:4982:151  */
  assign risone_d13 = n402; // (signal)
  /* fppow16.vhdl:4982:163  */
  assign risone_d14 = n403; // (signal)
  /* fppow16.vhdl:4982:175  */
  assign risone_d15 = n404; // (signal)
  /* fppow16.vhdl:4982:187  */
  assign risone_d16 = n405; // (signal)
  /* fppow16.vhdl:4982:199  */
  assign risone_d17 = n406; // (signal)
  /* fppow16.vhdl:4982:211  */
  assign risone_d18 = n407; // (signal)
  /* fppow16.vhdl:4982:223  */
  assign risone_d19 = n408; // (signal)
  /* fppow16.vhdl:4984:8  */
  assign risnan = n282; // (signal)
  /* fppow16.vhdl:4984:16  */
  assign risnan_d1 = n409; // (signal)
  /* fppow16.vhdl:4984:27  */
  assign risnan_d2 = n410; // (signal)
  /* fppow16.vhdl:4984:38  */
  assign risnan_d3 = n411; // (signal)
  /* fppow16.vhdl:4984:49  */
  assign risnan_d4 = n412; // (signal)
  /* fppow16.vhdl:4984:60  */
  assign risnan_d5 = n413; // (signal)
  /* fppow16.vhdl:4984:71  */
  assign risnan_d6 = n414; // (signal)
  /* fppow16.vhdl:4984:82  */
  assign risnan_d7 = n415; // (signal)
  /* fppow16.vhdl:4984:93  */
  assign risnan_d8 = n416; // (signal)
  /* fppow16.vhdl:4984:104  */
  assign risnan_d9 = n417; // (signal)
  /* fppow16.vhdl:4984:115  */
  assign risnan_d10 = n418; // (signal)
  /* fppow16.vhdl:4984:127  */
  assign risnan_d11 = n419; // (signal)
  /* fppow16.vhdl:4984:139  */
  assign risnan_d12 = n420; // (signal)
  /* fppow16.vhdl:4984:151  */
  assign risnan_d13 = n421; // (signal)
  /* fppow16.vhdl:4984:163  */
  assign risnan_d14 = n422; // (signal)
  /* fppow16.vhdl:4984:175  */
  assign risnan_d15 = n423; // (signal)
  /* fppow16.vhdl:4984:187  */
  assign risnan_d16 = n424; // (signal)
  /* fppow16.vhdl:4984:199  */
  assign risnan_d17 = n425; // (signal)
  /* fppow16.vhdl:4986:8  */
  assign signr = n283; // (signal)
  /* fppow16.vhdl:4986:15  */
  assign signr_d1 = n426; // (signal)
  /* fppow16.vhdl:4986:25  */
  assign signr_d2 = n427; // (signal)
  /* fppow16.vhdl:4986:35  */
  assign signr_d3 = n428; // (signal)
  /* fppow16.vhdl:4986:45  */
  assign signr_d4 = n429; // (signal)
  /* fppow16.vhdl:4986:55  */
  assign signr_d5 = n430; // (signal)
  /* fppow16.vhdl:4986:65  */
  assign signr_d6 = n431; // (signal)
  /* fppow16.vhdl:4986:75  */
  assign signr_d7 = n432; // (signal)
  /* fppow16.vhdl:4986:85  */
  assign signr_d8 = n433; // (signal)
  /* fppow16.vhdl:4986:95  */
  assign signr_d9 = n434; // (signal)
  /* fppow16.vhdl:4986:105  */
  assign signr_d10 = n435; // (signal)
  /* fppow16.vhdl:4986:116  */
  assign signr_d11 = n436; // (signal)
  /* fppow16.vhdl:4986:127  */
  assign signr_d12 = n437; // (signal)
  /* fppow16.vhdl:4986:138  */
  assign signr_d13 = n438; // (signal)
  /* fppow16.vhdl:4986:149  */
  assign signr_d14 = n439; // (signal)
  /* fppow16.vhdl:4986:160  */
  assign signr_d15 = n440; // (signal)
  /* fppow16.vhdl:4986:171  */
  assign signr_d16 = n441; // (signal)
  /* fppow16.vhdl:4986:182  */
  assign signr_d17 = n442; // (signal)
  /* fppow16.vhdl:4988:8  */
  assign login = n289; // (signal)
  /* fppow16.vhdl:4990:8  */
  assign lnx = fppow_5_10_freq500_uid2log_n290; // (signal)
  /* fppow16.vhdl:4992:8  */
  assign p = fppow_5_10_freq500_uid2mult_n293; // (signal)
  /* fppow16.vhdl:4994:8  */
  assign e = fppow_5_10_freq500_uid2exp_n296; // (signal)
  /* fppow16.vhdl:4994:11  */
  assign e_d1 = n443; // (signal)
  /* fppow16.vhdl:4996:8  */
  assign flagse = n299; // (signal)
  /* fppow16.vhdl:4996:16  */
  assign flagse_d1 = n444; // (signal)
  /* fppow16.vhdl:4998:8  */
  assign riszerofromexp = n303; // (signal)
  /* fppow16.vhdl:5000:8  */
  assign riszero = n305; // (signal)
  /* fppow16.vhdl:5002:8  */
  assign risinffromexp = n309; // (signal)
  /* fppow16.vhdl:5004:8  */
  assign risinf = n311; // (signal)
  /* fppow16.vhdl:5006:8  */
  assign flagr = n313; // (signal)
  /* fppow16.vhdl:5008:8  */
  assign r_expfrac = n320; // (signal)
  /* fppow16.vhdl:5139:15  */
  assign n126 = X[17:16]; // extract
  /* fppow16.vhdl:5140:14  */
  assign n127 = X[15]; // extract
  /* fppow16.vhdl:5141:18  */
  assign n128 = X[14:10]; // extract
  /* fppow16.vhdl:5142:14  */
  assign n129 = X[9:0]; // extract
  /* fppow16.vhdl:5143:15  */
  assign n130 = Y[17:16]; // extract
  /* fppow16.vhdl:5144:14  */
  assign n131 = Y[15]; // extract
  /* fppow16.vhdl:5145:18  */
  assign n132 = Y[14:10]; // extract
  /* fppow16.vhdl:5146:14  */
  assign n133 = Y[9:0]; // extract
  /* fppow16.vhdl:5149:28  */
  assign n136 = flagsx == 2'b00;
  /* fppow16.vhdl:5149:17  */
  assign n137 = n136 ? 1'b1 : 1'b0;
  /* fppow16.vhdl:5150:28  */
  assign n141 = flagsy == 2'b00;
  /* fppow16.vhdl:5150:17  */
  assign n142 = n141 ? 1'b1 : 1'b0;
  /* fppow16.vhdl:5152:30  */
  assign n146 = flagsx == 2'b01;
  /* fppow16.vhdl:5152:19  */
  assign n147 = n146 ? 1'b1 : 1'b0;
  /* fppow16.vhdl:5153:30  */
  assign n151 = flagsy == 2'b01;
  /* fppow16.vhdl:5153:19  */
  assign n152 = n151 ? 1'b1 : 1'b0;
  /* fppow16.vhdl:5155:27  */
  assign n156 = flagsx == 2'b10;
  /* fppow16.vhdl:5155:16  */
  assign n157 = n156 ? 1'b1 : 1'b0;
  /* fppow16.vhdl:5156:27  */
  assign n161 = flagsy == 2'b10;
  /* fppow16.vhdl:5156:16  */
  assign n162 = n161 ? 1'b1 : 1'b0;
  /* fppow16.vhdl:5158:31  */
  assign n166 = flagsx == 2'b11;
  /* fppow16.vhdl:5158:46  */
  assign n168 = flagsy == 2'b11;
  /* fppow16.vhdl:5158:37  */
  assign n169 = n166 | n168;
  /* fppow16.vhdl:5158:20  */
  assign n170 = n169 ? 1'b1 : 1'b0;
  /* fppow16.vhdl:5161:19  */
  assign n174 = {1'b0, expfieldx};
  /* fppow16.vhdl:5161:31  */
  assign n175 = {n174, fracx};
  /* fppow16.vhdl:5162:30  */
  assign n176 = ~oneexpfrac;
  /* fppow16.vhdl:5162:27  */
  assign n178 = {1'b1, n176};
  /* fppow16.vhdl:5163:4  */
  intadder_16_freq500_uid5 cmpxone (
    .clk(clk),
    .x(expfracx),
    .y(oneexpfraccompl),
    .cin(n179),
    .r(cmpxone_n180));
  /* fppow16.vhdl:5169:43  */
  assign n185 = {3'b010, oneexpfrac};
  /* fppow16.vhdl:5169:34  */
  assign n186 = X == n185;
  /* fppow16.vhdl:5169:27  */
  assign n187 = n186 ? 1'b1 : 1'b0;
  /* fppow16.vhdl:5170:39  */
  assign n189 = ~xisoneandnormal;
  /* fppow16.vhdl:5170:34  */
  assign n190 = normalx & n189;
  /* fppow16.vhdl:5170:79  */
  assign n191 = cmpxoneres[15]; // extract
  /* fppow16.vhdl:5170:65  */
  assign n192 = ~n191;
  /* fppow16.vhdl:5170:60  */
  assign n193 = n190 & n192;
  /* fppow16.vhdl:5171:48  */
  assign n194 = cmpxoneres[15]; // extract
  /* fppow16.vhdl:5171:34  */
  assign n195 = normalx & n194;
  /* fppow16.vhdl:5172:26  */
  assign n196 = fracy[0]; // extract
  /* fppow16.vhdl:5172:35  */
  assign n197 = fracy[1]; // extract
  /* fppow16.vhdl:5172:29  */
  assign n198 = {n196, n197};
  /* fppow16.vhdl:5172:44  */
  assign n199 = fracy[2]; // extract
  /* fppow16.vhdl:5172:38  */
  assign n200 = {n198, n199};
  /* fppow16.vhdl:5172:53  */
  assign n201 = fracy[3]; // extract
  /* fppow16.vhdl:5172:47  */
  assign n202 = {n200, n201};
  /* fppow16.vhdl:5172:62  */
  assign n203 = fracy[4]; // extract
  /* fppow16.vhdl:5172:56  */
  assign n204 = {n202, n203};
  /* fppow16.vhdl:5172:71  */
  assign n205 = fracy[5]; // extract
  /* fppow16.vhdl:5172:65  */
  assign n206 = {n204, n205};
  /* fppow16.vhdl:5172:80  */
  assign n207 = fracy[6]; // extract
  /* fppow16.vhdl:5172:74  */
  assign n208 = {n206, n207};
  /* fppow16.vhdl:5172:89  */
  assign n209 = fracy[7]; // extract
  /* fppow16.vhdl:5172:83  */
  assign n210 = {n208, n209};
  /* fppow16.vhdl:5172:98  */
  assign n211 = fracy[8]; // extract
  /* fppow16.vhdl:5172:92  */
  assign n212 = {n210, n211};
  /* fppow16.vhdl:5172:107  */
  assign n213 = fracy[9]; // extract
  /* fppow16.vhdl:5172:101  */
  assign n214 = {n212, n213};
  /* fppow16.vhdl:5173:4  */
  lzc_10_freq500_uid7 fppow_5_10_freq500_uid2right1counter (
    .clk(clk),
    .i(fracyreverted),
    .o(fppow_5_10_freq500_uid2right1counter_n215));
  /* fppow16.vhdl:5178:26  */
  assign n219 = {1'b0, expfieldy};
  /* fppow16.vhdl:5178:38  */
  assign n221 = n219 - 6'b011001;
  /* fppow16.vhdl:5179:35  */
  assign n222 = {2'b0, z_righty_d1};  //  uext
  /* fppow16.vhdl:5179:35  */
  assign n223 = weightlsbypre_d2 + n222;
  /* fppow16.vhdl:5180:42  */
  assign n225 = weightlsby == 6'b000000;
  /* fppow16.vhdl:5180:26  */
  assign n226 = n225 ? normaly_d2 : 1'b0;
  /* fppow16.vhdl:5181:42  */
  assign n228 = weightlsby[5]; // extract
  /* fppow16.vhdl:5181:46  */
  assign n229 = ~n228;
  /* fppow16.vhdl:5181:62  */
  assign n230 = ~oddinty;
  /* fppow16.vhdl:5181:51  */
  assign n231 = n230 & n229;
  /* fppow16.vhdl:5181:27  */
  assign n232 = n231 ? normaly_d2 : 1'b0;
  /* fppow16.vhdl:5182:47  */
  assign n234 = weightlsby[5]; // extract
  /* fppow16.vhdl:5182:32  */
  assign n235 = n234 ? normaly_d2 : 1'b0;
  /* fppow16.vhdl:5186:38  */
  assign n237 = oddinty_d1 | eveninty_d1;
  /* fppow16.vhdl:5186:21  */
  assign n238 = zerox_d3 & n237;
  /* fppow16.vhdl:5186:55  */
  assign n239 = n238 & signy_d3;
  /* fppow16.vhdl:5187:20  */
  assign n240 = zerox_d3 & infy_d3;
  /* fppow16.vhdl:5187:32  */
  assign n241 = n240 & signy_d3;
  /* fppow16.vhdl:5187:7  */
  assign n242 = n239 | n241;
  /* fppow16.vhdl:5188:35  */
  assign n243 = absxgtoneandnormal_d3 & infy_d3;
  /* fppow16.vhdl:5188:53  */
  assign n244 = ~signy_d3;
  /* fppow16.vhdl:5188:49  */
  assign n245 = n243 & n244;
  /* fppow16.vhdl:5188:7  */
  assign n246 = n242 | n245;
  /* fppow16.vhdl:5189:35  */
  assign n247 = absxltoneandnormal_d3 & infy_d3;
  /* fppow16.vhdl:5189:49  */
  assign n248 = n247 & signy_d3;
  /* fppow16.vhdl:5189:7  */
  assign n249 = n246 | n248;
  /* fppow16.vhdl:5190:19  */
  assign n250 = infx_d3 & normaly_d3;
  /* fppow16.vhdl:5190:40  */
  assign n251 = ~signy_d3;
  /* fppow16.vhdl:5190:36  */
  assign n252 = n250 & n251;
  /* fppow16.vhdl:5190:7  */
  assign n253 = n249 | n252;
  /* fppow16.vhdl:5192:37  */
  assign n254 = oddinty_d1 | eveninty_d1;
  /* fppow16.vhdl:5192:20  */
  assign n255 = zerox_d3 & n254;
  /* fppow16.vhdl:5192:58  */
  assign n256 = ~signy_d3;
  /* fppow16.vhdl:5192:54  */
  assign n257 = n255 & n256;
  /* fppow16.vhdl:5193:20  */
  assign n258 = zerox_d3 & infy_d3;
  /* fppow16.vhdl:5193:38  */
  assign n259 = ~signy_d3;
  /* fppow16.vhdl:5193:34  */
  assign n260 = n258 & n259;
  /* fppow16.vhdl:5193:7  */
  assign n261 = n257 | n260;
  /* fppow16.vhdl:5194:35  */
  assign n262 = absxltoneandnormal_d3 & infy_d3;
  /* fppow16.vhdl:5194:53  */
  assign n263 = ~signy_d3;
  /* fppow16.vhdl:5194:49  */
  assign n264 = n262 & n263;
  /* fppow16.vhdl:5194:7  */
  assign n265 = n261 | n264;
  /* fppow16.vhdl:5195:35  */
  assign n266 = absxgtoneandnormal_d3 & infy_d3;
  /* fppow16.vhdl:5195:49  */
  assign n267 = n266 & signy_d3;
  /* fppow16.vhdl:5195:7  */
  assign n268 = n265 | n267;
  /* fppow16.vhdl:5196:19  */
  assign n269 = infx_d3 & normaly_d3;
  /* fppow16.vhdl:5196:36  */
  assign n270 = n269 & signy_d3;
  /* fppow16.vhdl:5196:7  */
  assign n271 = n268 | n270;
  /* fppow16.vhdl:5199:27  */
  assign n272 = xisoneandnormal & signx;
  /* fppow16.vhdl:5199:37  */
  assign n273 = n272 & infy;
  /* fppow16.vhdl:5199:7  */
  assign n274 = zeroy | n273;
  /* fppow16.vhdl:5200:32  */
  assign n275 = ~signx;
  /* fppow16.vhdl:5200:28  */
  assign n276 = xisoneandnormal & n275;
  /* fppow16.vhdl:5200:7  */
  assign n277 = n274 | n276;
  /* fppow16.vhdl:5201:31  */
  assign n278 = ~zeroy_d2;
  /* fppow16.vhdl:5201:27  */
  assign n279 = s_nan_in_d2 & n278;
  /* fppow16.vhdl:5201:60  */
  assign n280 = normalx_d2 & signx_d2;
  /* fppow16.vhdl:5201:73  */
  assign n281 = n280 & notintnormaly;
  /* fppow16.vhdl:5201:45  */
  assign n282 = n279 | n281;
  /* fppow16.vhdl:5202:22  */
  assign n283 = signx_d2 & oddinty;
  /* fppow16.vhdl:5203:20  */
  assign n285 = {flagsx, 1'b0};
  /* fppow16.vhdl:5203:26  */
  assign n286 = {n285, expfieldx};
  /* fppow16.vhdl:5203:38  */
  assign n287 = {n286, fracx};
  /* fppow16.vhdl:5203:46  */
  assign n289 = {n287, 7'b0000000};
  /* fppow16.vhdl:5204:4  */
  fplogiterative_5_17_0_500_freq500_uid9 fppow_5_10_freq500_uid2log (
    .clk(clk),
    .x(login),
    .r(fppow_5_10_freq500_uid2log_n290));
  /* fppow16.vhdl:5208:4  */
  fpmult_5_17_uid57_freq500_uid58 fppow_5_10_freq500_uid2mult (
    .clk(clk),
    .x(lnx),
    .y(Y),
    .r(fppow_5_10_freq500_uid2mult_n293));
  /* fppow16.vhdl:5213:4  */
  fpexp_5_10_freq500_uid66 fppow_5_10_freq500_uid2exp (
    .clk(clk),
    .x(p),
    .r(fppow_5_10_freq500_uid2exp_n296));
  /* fppow16.vhdl:5217:15  */
  assign n299 = e[17:16]; // extract
  /* fppow16.vhdl:5218:40  */
  assign n302 = flagse_d1 == 2'b00;
  /* fppow16.vhdl:5218:26  */
  assign n303 = n302 ? 1'b1 : 1'b0;
  /* fppow16.vhdl:5219:38  */
  assign n305 = riszerospecialcase_d16 | riszerofromexp;
  /* fppow16.vhdl:5220:40  */
  assign n308 = flagse_d1 == 2'b10;
  /* fppow16.vhdl:5220:26  */
  assign n309 = n308 ? 1'b1 : 1'b0;
  /* fppow16.vhdl:5221:37  */
  assign n311 = risinfspecialcase_d16 | risinffromexp;
  /* fppow16.vhdl:5223:17  */
  assign n313 = risnan_d17 ? 2'b11 : n315;
  /* fppow16.vhdl:5224:7  */
  assign n315 = riszero ? 2'b00 : n317;
  /* fppow16.vhdl:5225:7  */
  assign n317 = risinf ? 2'b10 : 2'b01;
  /* fppow16.vhdl:5227:77  */
  assign n320 = risone_d19 ? 15'b011110000000000 : n321;
  /* fppow16.vhdl:5228:17  */
  assign n321 = e_d1[14:0]; // extract
  /* fppow16.vhdl:5229:15  */
  assign n322 = {flagr, signr_d17};
  /* fppow16.vhdl:5229:27  */
  assign n323 = {n322, r_expfrac};
  /* fppow16.vhdl:5015:10  */
  always @(posedge clk)
    n324 <= signx;
  /* fppow16.vhdl:5015:10  */
  always @(posedge clk)
    n325 <= signx_d1;
  /* fppow16.vhdl:5015:10  */
  always @(posedge clk)
    n326 <= signy;
  /* fppow16.vhdl:5015:10  */
  always @(posedge clk)
    n327 <= signy_d1;
  /* fppow16.vhdl:5015:10  */
  always @(posedge clk)
    n328 <= signy_d2;
  /* fppow16.vhdl:5015:10  */
  always @(posedge clk)
    n329 <= zerox;
  /* fppow16.vhdl:5015:10  */
  always @(posedge clk)
    n330 <= zerox_d1;
  /* fppow16.vhdl:5015:10  */
  always @(posedge clk)
    n331 <= zerox_d2;
  /* fppow16.vhdl:5015:10  */
  always @(posedge clk)
    n332 <= zeroy;
  /* fppow16.vhdl:5015:10  */
  always @(posedge clk)
    n333 <= zeroy_d1;
  /* fppow16.vhdl:5015:10  */
  always @(posedge clk)
    n334 <= normalx;
  /* fppow16.vhdl:5015:10  */
  always @(posedge clk)
    n335 <= normalx_d1;
  /* fppow16.vhdl:5015:10  */
  always @(posedge clk)
    n336 <= normaly;
  /* fppow16.vhdl:5015:10  */
  always @(posedge clk)
    n337 <= normaly_d1;
  /* fppow16.vhdl:5015:10  */
  always @(posedge clk)
    n338 <= normaly_d2;
  /* fppow16.vhdl:5015:10  */
  always @(posedge clk)
    n339 <= infx;
  /* fppow16.vhdl:5015:10  */
  always @(posedge clk)
    n340 <= infx_d1;
  /* fppow16.vhdl:5015:10  */
  always @(posedge clk)
    n341 <= infx_d2;
  /* fppow16.vhdl:5015:10  */
  always @(posedge clk)
    n342 <= infy;
  /* fppow16.vhdl:5015:10  */
  always @(posedge clk)
    n343 <= infy_d1;
  /* fppow16.vhdl:5015:10  */
  always @(posedge clk)
    n344 <= infy_d2;
  /* fppow16.vhdl:5015:10  */
  always @(posedge clk)
    n345 <= s_nan_in;
  /* fppow16.vhdl:5015:10  */
  always @(posedge clk)
    n346 <= s_nan_in_d1;
  /* fppow16.vhdl:5015:10  */
  always @(posedge clk)
    n347 <= absxgtoneandnormal;
  /* fppow16.vhdl:5015:10  */
  always @(posedge clk)
    n348 <= absxgtoneandnormal_d1;
  /* fppow16.vhdl:5015:10  */
  always @(posedge clk)
    n349 <= absxgtoneandnormal_d2;
  /* fppow16.vhdl:5015:10  */
  always @(posedge clk)
    n350 <= absxltoneandnormal;
  /* fppow16.vhdl:5015:10  */
  always @(posedge clk)
    n351 <= absxltoneandnormal_d1;
  /* fppow16.vhdl:5015:10  */
  always @(posedge clk)
    n352 <= absxltoneandnormal_d2;
  /* fppow16.vhdl:5015:10  */
  always @(posedge clk)
    n353 <= z_righty;
  /* fppow16.vhdl:5015:10  */
  always @(posedge clk)
    n354 <= weightlsbypre;
  /* fppow16.vhdl:5015:10  */
  always @(posedge clk)
    n355 <= weightlsbypre_d1;
  /* fppow16.vhdl:5015:10  */
  always @(posedge clk)
    n356 <= oddinty;
  /* fppow16.vhdl:5015:10  */
  always @(posedge clk)
    n357 <= eveninty;
  /* fppow16.vhdl:5015:10  */
  always @(posedge clk)
    n358 <= risinfspecialcase;
  /* fppow16.vhdl:5015:10  */
  always @(posedge clk)
    n359 <= risinfspecialcase_d1;
  /* fppow16.vhdl:5015:10  */
  always @(posedge clk)
    n360 <= risinfspecialcase_d2;
  /* fppow16.vhdl:5015:10  */
  always @(posedge clk)
    n361 <= risinfspecialcase_d3;
  /* fppow16.vhdl:5015:10  */
  always @(posedge clk)
    n362 <= risinfspecialcase_d4;
  /* fppow16.vhdl:5015:10  */
  always @(posedge clk)
    n363 <= risinfspecialcase_d5;
  /* fppow16.vhdl:5015:10  */
  always @(posedge clk)
    n364 <= risinfspecialcase_d6;
  /* fppow16.vhdl:5015:10  */
  always @(posedge clk)
    n365 <= risinfspecialcase_d7;
  /* fppow16.vhdl:5015:10  */
  always @(posedge clk)
    n366 <= risinfspecialcase_d8;
  /* fppow16.vhdl:5015:10  */
  always @(posedge clk)
    n367 <= risinfspecialcase_d9;
  /* fppow16.vhdl:5015:10  */
  always @(posedge clk)
    n368 <= risinfspecialcase_d10;
  /* fppow16.vhdl:5015:10  */
  always @(posedge clk)
    n369 <= risinfspecialcase_d11;
  /* fppow16.vhdl:5015:10  */
  always @(posedge clk)
    n370 <= risinfspecialcase_d12;
  /* fppow16.vhdl:5015:10  */
  always @(posedge clk)
    n371 <= risinfspecialcase_d13;
  /* fppow16.vhdl:5015:10  */
  always @(posedge clk)
    n372 <= risinfspecialcase_d14;
  /* fppow16.vhdl:5015:10  */
  always @(posedge clk)
    n373 <= risinfspecialcase_d15;
  /* fppow16.vhdl:5015:10  */
  always @(posedge clk)
    n374 <= riszerospecialcase;
  /* fppow16.vhdl:5015:10  */
  always @(posedge clk)
    n375 <= riszerospecialcase_d1;
  /* fppow16.vhdl:5015:10  */
  always @(posedge clk)
    n376 <= riszerospecialcase_d2;
  /* fppow16.vhdl:5015:10  */
  always @(posedge clk)
    n377 <= riszerospecialcase_d3;
  /* fppow16.vhdl:5015:10  */
  always @(posedge clk)
    n378 <= riszerospecialcase_d4;
  /* fppow16.vhdl:5015:10  */
  always @(posedge clk)
    n379 <= riszerospecialcase_d5;
  /* fppow16.vhdl:5015:10  */
  always @(posedge clk)
    n380 <= riszerospecialcase_d6;
  /* fppow16.vhdl:5015:10  */
  always @(posedge clk)
    n381 <= riszerospecialcase_d7;
  /* fppow16.vhdl:5015:10  */
  always @(posedge clk)
    n382 <= riszerospecialcase_d8;
  /* fppow16.vhdl:5015:10  */
  always @(posedge clk)
    n383 <= riszerospecialcase_d9;
  /* fppow16.vhdl:5015:10  */
  always @(posedge clk)
    n384 <= riszerospecialcase_d10;
  /* fppow16.vhdl:5015:10  */
  always @(posedge clk)
    n385 <= riszerospecialcase_d11;
  /* fppow16.vhdl:5015:10  */
  always @(posedge clk)
    n386 <= riszerospecialcase_d12;
  /* fppow16.vhdl:5015:10  */
  always @(posedge clk)
    n387 <= riszerospecialcase_d13;
  /* fppow16.vhdl:5015:10  */
  always @(posedge clk)
    n388 <= riszerospecialcase_d14;
  /* fppow16.vhdl:5015:10  */
  always @(posedge clk)
    n389 <= riszerospecialcase_d15;
  /* fppow16.vhdl:5015:10  */
  always @(posedge clk)
    n390 <= risone;
  /* fppow16.vhdl:5015:10  */
  always @(posedge clk)
    n391 <= risone_d1;
  /* fppow16.vhdl:5015:10  */
  always @(posedge clk)
    n392 <= risone_d2;
  /* fppow16.vhdl:5015:10  */
  always @(posedge clk)
    n393 <= risone_d3;
  /* fppow16.vhdl:5015:10  */
  always @(posedge clk)
    n394 <= risone_d4;
  /* fppow16.vhdl:5015:10  */
  always @(posedge clk)
    n395 <= risone_d5;
  /* fppow16.vhdl:5015:10  */
  always @(posedge clk)
    n396 <= risone_d6;
  /* fppow16.vhdl:5015:10  */
  always @(posedge clk)
    n397 <= risone_d7;
  /* fppow16.vhdl:5015:10  */
  always @(posedge clk)
    n398 <= risone_d8;
  /* fppow16.vhdl:5015:10  */
  always @(posedge clk)
    n399 <= risone_d9;
  /* fppow16.vhdl:5015:10  */
  always @(posedge clk)
    n400 <= risone_d10;
  /* fppow16.vhdl:5015:10  */
  always @(posedge clk)
    n401 <= risone_d11;
  /* fppow16.vhdl:5015:10  */
  always @(posedge clk)
    n402 <= risone_d12;
  /* fppow16.vhdl:5015:10  */
  always @(posedge clk)
    n403 <= risone_d13;
  /* fppow16.vhdl:5015:10  */
  always @(posedge clk)
    n404 <= risone_d14;
  /* fppow16.vhdl:5015:10  */
  always @(posedge clk)
    n405 <= risone_d15;
  /* fppow16.vhdl:5015:10  */
  always @(posedge clk)
    n406 <= risone_d16;
  /* fppow16.vhdl:5015:10  */
  always @(posedge clk)
    n407 <= risone_d17;
  /* fppow16.vhdl:5015:10  */
  always @(posedge clk)
    n408 <= risone_d18;
  /* fppow16.vhdl:5015:10  */
  always @(posedge clk)
    n409 <= risnan;
  /* fppow16.vhdl:5015:10  */
  always @(posedge clk)
    n410 <= risnan_d1;
  /* fppow16.vhdl:5015:10  */
  always @(posedge clk)
    n411 <= risnan_d2;
  /* fppow16.vhdl:5015:10  */
  always @(posedge clk)
    n412 <= risnan_d3;
  /* fppow16.vhdl:5015:10  */
  always @(posedge clk)
    n413 <= risnan_d4;
  /* fppow16.vhdl:5015:10  */
  always @(posedge clk)
    n414 <= risnan_d5;
  /* fppow16.vhdl:5015:10  */
  always @(posedge clk)
    n415 <= risnan_d6;
  /* fppow16.vhdl:5015:10  */
  always @(posedge clk)
    n416 <= risnan_d7;
  /* fppow16.vhdl:5015:10  */
  always @(posedge clk)
    n417 <= risnan_d8;
  /* fppow16.vhdl:5015:10  */
  always @(posedge clk)
    n418 <= risnan_d9;
  /* fppow16.vhdl:5015:10  */
  always @(posedge clk)
    n419 <= risnan_d10;
  /* fppow16.vhdl:5015:10  */
  always @(posedge clk)
    n420 <= risnan_d11;
  /* fppow16.vhdl:5015:10  */
  always @(posedge clk)
    n421 <= risnan_d12;
  /* fppow16.vhdl:5015:10  */
  always @(posedge clk)
    n422 <= risnan_d13;
  /* fppow16.vhdl:5015:10  */
  always @(posedge clk)
    n423 <= risnan_d14;
  /* fppow16.vhdl:5015:10  */
  always @(posedge clk)
    n424 <= risnan_d15;
  /* fppow16.vhdl:5015:10  */
  always @(posedge clk)
    n425 <= risnan_d16;
  /* fppow16.vhdl:5015:10  */
  always @(posedge clk)
    n426 <= signr;
  /* fppow16.vhdl:5015:10  */
  always @(posedge clk)
    n427 <= signr_d1;
  /* fppow16.vhdl:5015:10  */
  always @(posedge clk)
    n428 <= signr_d2;
  /* fppow16.vhdl:5015:10  */
  always @(posedge clk)
    n429 <= signr_d3;
  /* fppow16.vhdl:5015:10  */
  always @(posedge clk)
    n430 <= signr_d4;
  /* fppow16.vhdl:5015:10  */
  always @(posedge clk)
    n431 <= signr_d5;
  /* fppow16.vhdl:5015:10  */
  always @(posedge clk)
    n432 <= signr_d6;
  /* fppow16.vhdl:5015:10  */
  always @(posedge clk)
    n433 <= signr_d7;
  /* fppow16.vhdl:5015:10  */
  always @(posedge clk)
    n434 <= signr_d8;
  /* fppow16.vhdl:5015:10  */
  always @(posedge clk)
    n435 <= signr_d9;
  /* fppow16.vhdl:5015:10  */
  always @(posedge clk)
    n436 <= signr_d10;
  /* fppow16.vhdl:5015:10  */
  always @(posedge clk)
    n437 <= signr_d11;
  /* fppow16.vhdl:5015:10  */
  always @(posedge clk)
    n438 <= signr_d12;
  /* fppow16.vhdl:5015:10  */
  always @(posedge clk)
    n439 <= signr_d13;
  /* fppow16.vhdl:5015:10  */
  always @(posedge clk)
    n440 <= signr_d14;
  /* fppow16.vhdl:5015:10  */
  always @(posedge clk)
    n441 <= signr_d15;
  /* fppow16.vhdl:5015:10  */
  always @(posedge clk)
    n442 <= signr_d16;
  /* fppow16.vhdl:5015:10  */
  always @(posedge clk)
    n443 <= e;
  /* fppow16.vhdl:5015:10  */
  always @(posedge clk)
    n444 <= flagse;
endmodule

