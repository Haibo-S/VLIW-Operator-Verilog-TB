--------------------------------------------------------------------------------
--                          InvA0Table_Freq500_uid15
-- VHDL generated for DummyFPGA @ 500MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 2
-- Target frequency (MHz): 500
-- Input signals: X
-- Output signals: Y
--  approx. input signal timings: X: (c0, 0.000000ns)
--  approx. output signal timings: Y: (c0, 0.550000ns)

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity InvA0Table_Freq500_uid15 is
    port (X : in  std_logic_vector(7 downto 0);
          Y : out  std_logic_vector(8 downto 0)   );
end entity;

architecture arch of InvA0Table_Freq500_uid15 is
signal Y0 :  std_logic_vector(8 downto 0);
   -- timing of Y0: (c0, 0.550000ns)
signal Y1 :  std_logic_vector(8 downto 0);
   -- timing of Y1: (c0, 0.550000ns)
begin
   with X  select  Y0 <= 
      "100000000" when "00000000",
      "100000000" when "00000001",
      "011111111" when "00000010",
      "011111110" when "00000011",
      "011111101" when "00000100",
      "011111100" when "00000101",
      "011111011" when "00000110",
      "011111010" when "00000111",
      "011111001" when "00001000",
      "011111000" when "00001001",
      "011110111" when "00001010",
      "011110110" when "00001011",
      "011110101" when "00001100",
      "011110100" when "00001101",
      "011110011" when "00001110",
      "011110010" when "00001111",
      "011110001" when "00010000",
      "011110001" when "00010001",
      "011110000" when "00010010",
      "011101111" when "00010011",
      "011101110" when "00010100",
      "011101101" when "00010101",
      "011101100" when "00010110",
      "011101011" when "00010111",
      "011101011" when "00011000",
      "011101010" when "00011001",
      "011101001" when "00011010",
      "011101000" when "00011011",
      "011100111" when "00011100",
      "011100110" when "00011101",
      "011100110" when "00011110",
      "011100101" when "00011111",
      "011100100" when "00100000",
      "011100011" when "00100001",
      "011100010" when "00100010",
      "011100010" when "00100011",
      "011100001" when "00100100",
      "011100000" when "00100101",
      "011011111" when "00100110",
      "011011111" when "00100111",
      "011011110" when "00101000",
      "011011101" when "00101001",
      "011011100" when "00101010",
      "011011100" when "00101011",
      "011011011" when "00101100",
      "011011010" when "00101101",
      "011011010" when "00101110",
      "011011001" when "00101111",
      "011011000" when "00110000",
      "011010111" when "00110001",
      "011010111" when "00110010",
      "011010110" when "00110011",
      "011010101" when "00110100",
      "011010101" when "00110101",
      "011010100" when "00110110",
      "011010011" when "00110111",
      "011010011" when "00111000",
      "011010010" when "00111001",
      "011010001" when "00111010",
      "011010001" when "00111011",
      "011010000" when "00111100",
      "011001111" when "00111101",
      "011001111" when "00111110",
      "011001110" when "00111111",
      "011001101" when "01000000",
      "011001101" when "01000001",
      "011001100" when "01000010",
      "011001011" when "01000011",
      "011001011" when "01000100",
      "011001010" when "01000101",
      "011001010" when "01000110",
      "011001001" when "01000111",
      "011001000" when "01001000",
      "011001000" when "01001001",
      "011000111" when "01001010",
      "011000110" when "01001011",
      "011000110" when "01001100",
      "011000101" when "01001101",
      "011000101" when "01001110",
      "011000100" when "01001111",
      "011000100" when "01010000",
      "011000011" when "01010001",
      "011000010" when "01010010",
      "011000010" when "01010011",
      "011000001" when "01010100",
      "011000001" when "01010101",
      "011000000" when "01010110",
      "011000000" when "01010111",
      "010111111" when "01011000",
      "010111110" when "01011001",
      "010111110" when "01011010",
      "010111101" when "01011011",
      "010111101" when "01011100",
      "010111100" when "01011101",
      "010111100" when "01011110",
      "010111011" when "01011111",
      "010111011" when "01100000",
      "010111010" when "01100001",
      "010111010" when "01100010",
      "010111001" when "01100011",
      "010111001" when "01100100",
      "010111000" when "01100101",
      "010111000" when "01100110",
      "010110111" when "01100111",
      "010110111" when "01101000",
      "010110110" when "01101001",
      "010110110" when "01101010",
      "010110101" when "01101011",
      "010110101" when "01101100",
      "010110100" when "01101101",
      "010110100" when "01101110",
      "010110011" when "01101111",
      "010110011" when "01110000",
      "010110010" when "01110001",
      "010110010" when "01110010",
      "010110001" when "01110011",
      "010110001" when "01110100",
      "010110000" when "01110101",
      "010110000" when "01110110",
      "010101111" when "01110111",
      "010101111" when "01111000",
      "010101110" when "01111001",
      "010101110" when "01111010",
      "010101101" when "01111011",
      "010101101" when "01111100",
      "010101101" when "01111101",
      "010101100" when "01111110",
      "010101100" when "01111111",
      "101010110" when "10000000",
      "101010101" when "10000001",
      "101010100" when "10000010",
      "101010011" when "10000011",
      "101010010" when "10000100",
      "101010001" when "10000101",
      "101010001" when "10000110",
      "101010000" when "10000111",
      "101001111" when "10001000",
      "101001110" when "10001001",
      "101001101" when "10001010",
      "101001100" when "10001011",
      "101001011" when "10001100",
      "101001011" when "10001101",
      "101001010" when "10001110",
      "101001001" when "10001111",
      "101001000" when "10010000",
      "101000111" when "10010001",
      "101000111" when "10010010",
      "101000110" when "10010011",
      "101000101" when "10010100",
      "101000100" when "10010101",
      "101000011" when "10010110",
      "101000011" when "10010111",
      "101000010" when "10011000",
      "101000001" when "10011001",
      "101000000" when "10011010",
      "100111111" when "10011011",
      "100111111" when "10011100",
      "100111110" when "10011101",
      "100111101" when "10011110",
      "100111100" when "10011111",
      "100111100" when "10100000",
      "100111011" when "10100001",
      "100111010" when "10100010",
      "100111001" when "10100011",
      "100111001" when "10100100",
      "100111000" when "10100101",
      "100110111" when "10100110",
      "100110110" when "10100111",
      "100110110" when "10101000",
      "100110101" when "10101001",
      "100110100" when "10101010",
      "100110011" when "10101011",
      "100110011" when "10101100",
      "100110010" when "10101101",
      "100110001" when "10101110",
      "100110001" when "10101111",
      "100110000" when "10110000",
      "100101111" when "10110001",
      "100101111" when "10110010",
      "100101110" when "10110011",
      "100101101" when "10110100",
      "100101100" when "10110101",
      "100101100" when "10110110",
      "100101011" when "10110111",
      "100101010" when "10111000",
      "100101010" when "10111001",
      "100101001" when "10111010",
      "100101000" when "10111011",
      "100101000" when "10111100",
      "100100111" when "10111101",
      "100100110" when "10111110",
      "100100110" when "10111111",
      "100100101" when "11000000",
      "100100100" when "11000001",
      "100100100" when "11000010",
      "100100011" when "11000011",
      "100100010" when "11000100",
      "100100010" when "11000101",
      "100100001" when "11000110",
      "100100001" when "11000111",
      "100100000" when "11001000",
      "100011111" when "11001001",
      "100011111" when "11001010",
      "100011110" when "11001011",
      "100011101" when "11001100",
      "100011101" when "11001101",
      "100011100" when "11001110",
      "100011100" when "11001111",
      "100011011" when "11010000",
      "100011010" when "11010001",
      "100011010" when "11010010",
      "100011001" when "11010011",
      "100011001" when "11010100",
      "100011000" when "11010101",
      "100010111" when "11010110",
      "100010111" when "11010111",
      "100010110" when "11011000",
      "100010110" when "11011001",
      "100010101" when "11011010",
      "100010100" when "11011011",
      "100010100" when "11011100",
      "100010011" when "11011101",
      "100010011" when "11011110",
      "100010010" when "11011111",
      "100010010" when "11100000",
      "100010001" when "11100001",
      "100010000" when "11100010",
      "100010000" when "11100011",
      "100001111" when "11100100",
      "100001111" when "11100101",
      "100001110" when "11100110",
      "100001110" when "11100111",
      "100001101" when "11101000",
      "100001101" when "11101001",
      "100001100" when "11101010",
      "100001011" when "11101011",
      "100001011" when "11101100",
      "100001010" when "11101101",
      "100001010" when "11101110",
      "100001001" when "11101111",
      "100001001" when "11110000",
      "100001000" when "11110001",
      "100001000" when "11110010",
      "100000111" when "11110011",
      "100000111" when "11110100",
      "100000110" when "11110101",
      "100000110" when "11110110",
      "100000101" when "11110111",
      "100000101" when "11111000",
      "100000100" when "11111001",
      "100000100" when "11111010",
      "100000011" when "11111011",
      "100000011" when "11111100",
      "100000010" when "11111101",
      "100000010" when "11111110",
      "100000001" when "11111111",
      "---------" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          LogTable0_Freq500_uid27
-- VHDL generated for DummyFPGA @ 500MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 2
-- Target frequency (MHz): 500
-- Input signals: X
-- Output signals: Y
--  approx. input signal timings: X: (c0, 0.000000ns)
--  approx. output signal timings: Y: (c0, 0.550000ns)

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity LogTable0_Freq500_uid27 is
    port (X : in  std_logic_vector(7 downto 0);
          Y : out  std_logic_vector(34 downto 0)   );
end entity;

architecture arch of LogTable0_Freq500_uid27 is
signal Y0 :  std_logic_vector(34 downto 0);
   -- timing of Y0: (c0, 0.550000ns)
signal Y1 :  std_logic_vector(34 downto 0);
   -- timing of Y1: (c0, 0.550000ns)
begin
   with X  select  Y0 <= 
      "11111111111100000000000000000000000" when "00000000",
      "11111111111100000000000000000000000" when "00000001",
      "00000000111100001000000001010101101" when "00000010",
      "00000001111100100000001010101110110" when "00000011",
      "00000010111101001000100100010100100" when "00000100",
      "00000011111110000001010110010110001" when "00000101",
      "00000100111111001010101001001001011" when "00000110",
      "00000110000000100100100101001010010" when "00000111",
      "00000111000010001111010010111011000" when "00001000",
      "00001000000100001010111011000101000" when "00001001",
      "00001001000110010111100110010111110" when "00001010",
      "00001010001000110101011101101010001" when "00001011",
      "00001011001011100100101001111001011" when "00001100",
      "00001100001110100101010100001010010" when "00001101",
      "00001101010001110111100101101000100" when "00001110",
      "00001110010101011011100111100110111" when "00001111",
      "00001111011001010001100011100000000" when "00010000",
      "00001111011001010001100011100000000" when "00010001",
      "00010000011101011001100010110101101" when "00010010",
      "00010001100001110011101111010001010" when "00010011",
      "00010010100110100000010010100100010" when "00010100",
      "00010011101011011111010110100111110" when "00010101",
      "00010100110000110001000101011101001" when "00010110",
      "00010101110110010101101001001101101" when "00010111",
      "00010101110110010101101001001101101" when "00011000",
      "00010110111100001101001100001010111" when "00011001",
      "00011000000010010111111000101111010" when "00011010",
      "00011001001000110101111001011101011" when "00011011",
      "00011010001111100111011001000000110" when "00011100",
      "00011011010110101100100010001101101" when "00011101",
      "00011011010110101100100010001101101" when "00011110",
      "00011100011110000101100000000001110" when "00011111",
      "00011101100101110010011101100011100" when "00100000",
      "00011110101101110011100110000011000" when "00100001",
      "00011111110110001001000100111001111" when "00100010",
      "00011111110110001001000100111001111" when "00100011",
      "00100000111110110011000101101011010" when "00100100",
      "00100010000111110001110100000100010" when "00100101",
      "00100011010001000101011011111100010" when "00100110",
      "00100011010001000101011011111100010" when "00100111",
      "00100100011010101110001001010100100" when "00101000",
      "00100101100100101100001000011001000" when "00101001",
      "00100110101110111111100101100000001" when "00101010",
      "00100110101110111111100101100000001" when "00101011",
      "00100111111001101000101101001011010" when "00101100",
      "00101001000100100111101100000110011" when "00101101",
      "00101001000100100111101100000110011" when "00101110",
      "00101010001111111100101111001001010" when "00101111",
      "00101011011011101000000011010110101" when "00110000",
      "00101100100111101001110101111101001" when "00110001",
      "00101100100111101001110101111101001" when "00110010",
      "00101101110100000010010100010110111" when "00110011",
      "00101111000000110001101100001010100" when "00110100",
      "00101111000000110001101100001010100" when "00110101",
      "00110000001101111000001011001010101" when "00110110",
      "00110001011011010101111111010110100" when "00110111",
      "00110001011011010101111111010110100" when "00111000",
      "00110010101001001011010110111010000" when "00111001",
      "00110011110111011000100000001110000" when "00111010",
      "00110011110111011000100000001110000" when "00111011",
      "00110101000101111101101001111001001" when "00111100",
      "00110110010100111011000010101110110" when "00111101",
      "00110110010100111011000010101110110" when "00111110",
      "00110111100100010000111001110000100" when "00111111",
      "00111000110011111111011110001101111" when "01000000",
      "00111000110011111111011110001101111" when "01000001",
      "00111010000100000110111111100100110" when "01000010",
      "00111011010100100111101101100001101" when "01000011",
      "00111011010100100111101101100001101" when "01000100",
      "00111100100101100001110111111111110" when "01000101",
      "00111100100101100001110111111111110" when "01000110",
      "00111101110110110101101111001001110" when "01000111",
      "00111111001000100011100011011001011" when "01001000",
      "00111111001000100011100011011001011" when "01001001",
      "01000000011010101011100101011000101" when "01001010",
      "01000001101101001110000110000001010" when "01001011",
      "01000001101101001110000110000001010" when "01001100",
      "01000011000000001011010110011101100" when "01001101",
      "01000011000000001011010110011101100" when "01001110",
      "01000100010011100011101000001000101" when "01001111",
      "01000100010011100011101000001000101" when "01010000",
      "01000101100111010111001100101110110" when "01010001",
      "01000110111011100110010110001101100" when "01010010",
      "01000110111011100110010110001101100" when "01010011",
      "01001000010000010001010110110100010" when "01010100",
      "01001000010000010001010110110100010" when "01010101",
      "01001001100101011000100001000100110" when "01010110",
      "01001001100101011000100001000100110" when "01010111",
      "01001010111010111100000111110011100" when "01011000",
      "01001100010000111100011110000111010" when "01011001",
      "01001100010000111100011110000111010" when "01011010",
      "01001101100111011001110111011011000" when "01011011",
      "01001101100111011001110111011011000" when "01011100",
      "01001110111110010100100111011100110" when "01011101",
      "01001110111110010100100111011100110" when "01011110",
      "01010000010101101101000010001111010" when "01011111",
      "01010000010101101101000010001111010" when "01100000",
      "01010001101101100011011100001001110" when "01100001",
      "01010001101101100011011100001001110" when "01100010",
      "01010011000101111000001001111000011" when "01100011",
      "01010011000101111000001001111000011" when "01100100",
      "01010100011110101011100000011100111" when "01100101",
      "01010100011110101011100000011100111" when "01100110",
      "01010101110111111101110101001111001" when "01100111",
      "01010101110111111101110101001111001" when "01101000",
      "01010111010001101111011101111101011" when "01101001",
      "01010111010001101111011101111101011" when "01101010",
      "01011000101100000000110000101101000" when "01101011",
      "01011000101100000000110000101101000" when "01101100",
      "01011010000110110010000011111010100" when "01101101",
      "01011010000110110010000011111010100" when "01101110",
      "01011011100010000011101110011010110" when "01101111",
      "01011011100010000011101110011010110" when "01110000",
      "01011100111101110110000111011011001" when "01110001",
      "01011100111101110110000111011011001" when "01110010",
      "01011110011010001001100110100010000" when "01110011",
      "01011110011010001001100110100010000" when "01110100",
      "01011111110110111110100011101111011" when "01110101",
      "01011111110110111110100011101111011" when "01110110",
      "01100001010100010101010111011101110" when "01110111",
      "01100001010100010101010111011101110" when "01111000",
      "01100010110010001110011010100010010" when "01111001",
      "01100010110010001110011010100010010" when "01111010",
      "01100100010000101010000110001101100" when "01111011",
      "01100100010000101010000110001101100" when "01111100",
      "01100100010000101010000110001101100" when "01111101",
      "01100101101111101000110100001100010" when "01111110",
      "01100101101111101000110100001100010" when "01111111",
      "10110101110010101001011110110000100" when "10000000",
      "10110110100010100111111110111100100" when "10000001",
      "10110111010010101111100000010000110" when "10000010",
      "10111000000011000000000110000110111" when "10000011",
      "10111000110011011001110011111010011" when "10000100",
      "10111001100011111100101101001000110" when "10000101",
      "10111001100011111100101101001000110" when "10000110",
      "10111010010100101000110101010001010" when "10000111",
      "10111011000101011110001111110101110" when "10001000",
      "10111011110110011101000000011001010" when "10001001",
      "10111100100111100101001010100001100" when "10001010",
      "10111101011000110110110001110110010" when "10001011",
      "10111110001010010001111010000000110" when "10001100",
      "10111110001010010001111010000000110" when "10001101",
      "10111110111011110110100110101101010" when "10001110",
      "10111111101101100100111011101001010" when "10001111",
      "11000000011111011100111100100101010" when "10010000",
      "11000001010001011110101101010011011" when "10010001",
      "11000001010001011110101101010011011" when "10010010",
      "11000010000011101010010001101000010" when "10010011",
      "11000010110101111111101101011010101" when "10010100",
      "11000011101000011111000100100011101" when "10010101",
      "11000100011011001000011010111110101" when "10010110",
      "11000100011011001000011010111110101" when "10010111",
      "11000101001101111011110100101001011" when "10011000",
      "11000110000000111001010101100100000" when "10011001",
      "11000110110100000001000001110000110" when "10011010",
      "11000111100111010010111101010100111" when "10011011",
      "11000111100111010010111101010100111" when "10011100",
      "11001000011010101111001100010111101" when "10011101",
      "11001001001110010101110011000010111" when "10011110",
      "11001010000010000110110101100011000" when "10011111",
      "11001010000010000110110101100011000" when "10100000",
      "11001010110110000010011000000111000" when "10100001",
      "11001011101010001000011111000000010" when "10100010",
      "11001100011110011001001110100011000" when "10100011",
      "11001100011110011001001110100011000" when "10100100",
      "11001101010010110100101011000110001" when "10100101",
      "11001110000111011010111001000011000" when "10100110",
      "11001110111100001011111100110101110" when "10100111",
      "11001110111100001011111100110101110" when "10101000",
      "11001111110001000111111010111101100" when "10101001",
      "11010000100110001110110111111011111" when "10101010",
      "11010001011011100000111000010101100" when "10101011",
      "11010001011011100000111000010101100" when "10101100",
      "11010010010000111110000000110001110" when "10101101",
      "11010011000110100110010101111011001" when "10101110",
      "11010011000110100110010101111011001" when "10101111",
      "11010011111100011001111100011110110" when "10110000",
      "11010100110010011000111001001100110" when "10110001",
      "11010100110010011000111001001100110" when "10110010",
      "11010101101000100011010000111000110" when "10110011",
      "11010110011110111001001000011000110" when "10110100",
      "11010111010101011010100100100110011" when "10110101",
      "11010111010101011010100100100110011" when "10110110",
      "11011000001100000111101010011110001" when "10110111",
      "11011001000011000000011110111111110" when "10111000",
      "11011001000011000000011110111111110" when "10111001",
      "11011001111010000101000111001110010" when "10111010",
      "11011010110001010101101000001111110" when "10111011",
      "11011010110001010101101000001111110" when "10111100",
      "11011011101000110010000111001101111" when "10111101",
      "11011100100000011010101001010101101" when "10111110",
      "11011100100000011010101001010101101" when "10111111",
      "11011101011000001111010011110111010" when "11000000",
      "11011110010000010000001100000110011" when "11000001",
      "11011110010000010000001100000110011" when "11000010",
      "11011111001000011101010111011010011" when "11000011",
      "11100000000000110110111011001110001" when "11000100",
      "11100000000000110110111011001110001" when "11000101",
      "11100000111001011100111101000000000" when "11000110",
      "11100000111001011100111101000000000" when "11000111",
      "11100001110010001111100010010001111" when "11001000",
      "11100010101011001110110000101001101" when "11001001",
      "11100010101011001110110000101001101" when "11001010",
      "11100011100100011010101101110000101" when "11001011",
      "11100100011101110011011111010100010" when "11001100",
      "11100100011101110011011111010100010" when "11001101",
      "11100101010111011001001011000101110" when "11001110",
      "11100101010111011001001011000101110" when "11001111",
      "11100110010001001011110110111001111" when "11010000",
      "11100111001011001011101000101001110" when "11010001",
      "11100111001011001011101000101001110" when "11010010",
      "11101000000101011000100110010010100" when "11010011",
      "11101000000101011000100110010010100" when "11010100",
      "11101000111111110010110101110101001" when "11010101",
      "11101001111010011010011101010110110" when "11010110",
      "11101001111010011010011101010110110" when "11010111",
      "11101010110101001111100011000001000" when "11011000",
      "11101010110101001111100011000001000" when "11011001",
      "11101011110000010010001101000001011" when "11011010",
      "11101100101011100010100001101001111" when "11011011",
      "11101100101011100010100001101001111" when "11011100",
      "11101101100111000000100111010001000" when "11011101",
      "11101101100111000000100111010001000" when "11011110",
      "11101110100010101100100100010001011" when "11011111",
      "11101110100010101100100100010001011" when "11100000",
      "11101111011110100110011111001010011" when "11100001",
      "11110000011010101110011110100000000" when "11100010",
      "11110000011010101110011110100000000" when "11100011",
      "11110001010111000100101000111010101" when "11100100",
      "11110001010111000100101000111010101" when "11100101",
      "11110010010011101001000101000111100" when "11100110",
      "11110010010011101001000101000111100" when "11100111",
      "11110011010000011011111001111000101" when "11101000",
      "11110011010000011011111001111000101" when "11101001",
      "11110100001101011101001110000100111" when "11101010",
      "11110101001010101101001000101000001" when "11101011",
      "11110101001010101101001000101000001" when "11101100",
      "11110110001000001011110000100011000" when "11101101",
      "11110110001000001011110000100011000" when "11101110",
      "11110111000101111001001100111011011" when "11101111",
      "11110111000101111001001100111011011" when "11110000",
      "11111000000011110101100100111100011" when "11110001",
      "11111000000011110101100100111100011" when "11110010",
      "11111001000010000000111111110110001" when "11110011",
      "11111001000010000000111111110110001" when "11110100",
      "11111010000000011011100100111110000" when "11110101",
      "11111010000000011011100100111110000" when "11110110",
      "11111010111111000101011011101111001" when "11110111",
      "11111010111111000101011011101111001" when "11111000",
      "11111011111101111110101011101001111" when "11111001",
      "11111011111101111110101011101001111" when "11111010",
      "11111100111101000111011100010100000" when "11111011",
      "11111100111101000111011100010100000" when "11111100",
      "11111101111100011111110101011001010" when "11111101",
      "11111101111100011111110101011001010" when "11111110",
      "11111110111100000111111110101010111" when "11111111",
      "-----------------------------------" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          LogTable1_Freq500_uid30
-- VHDL generated for DummyFPGA @ 500MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 2
-- Target frequency (MHz): 500
-- Input signals: X
-- Output signals: Y
--  approx. input signal timings: X: (c0, 0.000000ns)
--  approx. output signal timings: Y: (c0, 0.600000ns)

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity LogTable1_Freq500_uid30 is
    port (X : in  std_logic_vector(5 downto 0);
          Y : out  std_logic_vector(28 downto 0)   );
end entity;

architecture arch of LogTable1_Freq500_uid30 is
signal Y0 :  std_logic_vector(28 downto 0);
   -- timing of Y0: (c0, 0.600000ns)
signal Y1 :  std_logic_vector(28 downto 0);
   -- timing of Y1: (c0, 0.600000ns)
begin
   with X  select  Y0 <= 
      "00000010000000000000100000000" when "000000",
      "00000110000000000000100000000" when "000001",
      "00001010000000000100100000001" when "000010",
      "00001110000000001100100000011" when "000011",
      "00010010000000011000100000111" when "000100",
      "00010110000000101000100001111" when "000101",
      "00011010000000111100100011100" when "000110",
      "00011110000001010100100101110" when "000111",
      "00100010000001110000101000110" when "001000",
      "00100110000010010000101100110" when "001001",
      "00101010000010110100110001111" when "001010",
      "00101110000011011100111000001" when "001011",
      "00110010000100001000111111110" when "001100",
      "00110110000100111001001000110" when "001101",
      "00111010000101101101010011011" when "001110",
      "00111110000110100101011111110" when "001111",
      "01000010000111100001101101110" when "010000",
      "01000110001000100001111101111" when "010001",
      "01001010001001100110010000000" when "010010",
      "01001110001010101110100100011" when "010011",
      "01010010001011111010111011000" when "010100",
      "01010110001101001011010100010" when "010101",
      "01011010001110011111101111111" when "010110",
      "01011110001111111000001110010" when "010111",
      "01100010010001010100101111100" when "011000",
      "01100110010010110101010011110" when "011001",
      "01101010010100011001111011000" when "011010",
      "01101110010110000010100101100" when "011011",
      "01110010010111101111010011100" when "011100",
      "01110110011001100000000100110" when "011101",
      "01111010011011010100111001110" when "011110",
      "01111110011101001101110010100" when "011111",
      "10000000011110001011110000010" when "100000",
      "10000100100000001010101110110" when "100001",
      "10001000100010001101110001010" when "100010",
      "10001100100100010100111000000" when "100011",
      "10010000100110100000000011000" when "100100",
      "10010100101000101111010010100" when "100101",
      "10011000101011000010100110100" when "100110",
      "10011100101101011001111111001" when "100111",
      "10100000101111110101011100110" when "101000",
      "10100100110010010100111111001" when "101001",
      "10101000110100111000100110110" when "101010",
      "10101100110111100000010011100" when "101011",
      "10110000111010001100000101100" when "101100",
      "10110100111100111011111101001" when "101101",
      "10111000111111101111111010010" when "101110",
      "10111101000010100111111101001" when "101111",
      "11000001000101100100000101110" when "110000",
      "11000101001000100100010100100" when "110001",
      "11001001001011101000101001010" when "110010",
      "11001101001110110001000100010" when "110011",
      "11010001010001111101100101101" when "110100",
      "11010101010101001110001101100" when "110101",
      "11011001011000100010111100000" when "110110",
      "11011101011011111011110001010" when "110111",
      "11100001011111011000101101011" when "111000",
      "11100101100010111001110000101" when "111001",
      "11101001100110011110111010111" when "111010",
      "11101101101010001000001100100" when "111011",
      "11110001101101110101100101100" when "111100",
      "11110101110001100111000110000" when "111101",
      "11111001110101011100101110010" when "111110",
      "11111101111001010110011110010" when "111111",
      "-----------------------------" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                 FixRealKCM_Freq500_uid39_T0_Freq500_uid42
-- VHDL generated for DummyFPGA @ 500MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 2
-- Target frequency (MHz): 500
-- Input signals: X
-- Output signals: Y
--  approx. input signal timings: X: (c0, 0.000000ns)
--  approx. output signal timings: Y: (c0, 0.550000ns)

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity FixRealKCM_Freq500_uid39_T0_Freq500_uid42 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(31 downto 0)   );
end entity;

architecture arch of FixRealKCM_Freq500_uid39_T0_Freq500_uid42 is
signal Y0 :  std_logic_vector(31 downto 0);
   -- timing of Y0: (c0, 0.550000ns)
signal Y1 :  std_logic_vector(31 downto 0);
   -- timing of Y1: (c0, 0.550000ns)
begin
   with X  select  Y0 <= 
      "00000000000000000000000000000000" when "00000",
      "00000101100010111001000011000000" when "00001",
      "00001011000101110010000101111111" when "00010",
      "00010000101000101011001000111111" when "00011",
      "00010110001011100100001011111111" when "00100",
      "00011011101110011101001110111111" when "00101",
      "00100001010001010110010001111110" when "00110",
      "00100110110100001111010100111110" when "00111",
      "00101100010111001000010111111110" when "01000",
      "00110001111010000001011010111110" when "01001",
      "00110111011100111010011101111101" when "01010",
      "00111100111111110011100000111101" when "01011",
      "01000010100010101100100011111101" when "01100",
      "01001000000101100101100110111101" when "01101",
      "01001101101000011110101001111100" when "01110",
      "01010011001011010111101100111100" when "01111",
      "01011000101110010000101111111100" when "10000",
      "01011110010001001001110010111100" when "10001",
      "01100011110100000010110101111011" when "10010",
      "01101001010110111011111000111011" when "10011",
      "01101110111001110100111011111011" when "10100",
      "01110100011100101101111110111011" when "10101",
      "01111001111111100111000001111010" when "10110",
      "01111111100010100000000100111010" when "10111",
      "10000101000101011001000111111010" when "11000",
      "10001010101000010010001010111010" when "11001",
      "10010000001011001011001101111001" when "11010",
      "10010101101110000100010000111001" when "11011",
      "10011011010000111101010011111001" when "11100",
      "10100000110011110110010110111001" when "11101",
      "10100110010110101111011001111000" when "11110",
      "10101011111001101000011100111000" when "11111",
      "--------------------------------" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                 FixRealKCM_Freq500_uid39_T1_Freq500_uid45
-- VHDL generated for DummyFPGA @ 500MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 2
-- Target frequency (MHz): 500
-- Input signals: X
-- Output signals: Y
--  approx. input signal timings: X: (c0, 0.000000ns)
--  approx. output signal timings: Y: (c0, 0.550000ns)

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity FixRealKCM_Freq500_uid39_T1_Freq500_uid45 is
    port (X : in  std_logic_vector(2 downto 0);
          Y : out  std_logic_vector(26 downto 0)   );
end entity;

architecture arch of FixRealKCM_Freq500_uid39_T1_Freq500_uid45 is
signal Y0 :  std_logic_vector(26 downto 0);
   -- timing of Y0: (c0, 0.550000ns)
signal Y1 :  std_logic_vector(26 downto 0);
   -- timing of Y1: (c0, 0.550000ns)
begin
   with X  select  Y0 <= 
      "000000000000000000000000000" when "000",
      "000101100010111001000011000" when "001",
      "001011000101110010000110000" when "010",
      "010000101000101011001001000" when "011",
      "010110001011100100001100000" when "100",
      "011011101110011101001111000" when "101",
      "100001010001010110010010000" when "110",
      "100110110100001111010101000" when "111",
      "---------------------------" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                 FixRealKCM_Freq500_uid77_T0_Freq500_uid80
-- VHDL generated for DummyFPGA @ 500MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 2
-- Target frequency (MHz): 500
-- Input signals: X
-- Output signals: Y
--  approx. input signal timings: X: (c0, 0.000000ns)
--  approx. output signal timings: Y: (c0, 0.550000ns)

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity FixRealKCM_Freq500_uid77_T0_Freq500_uid80 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(11 downto 0)   );
end entity;

architecture arch of FixRealKCM_Freq500_uid77_T0_Freq500_uid80 is
signal Y0 :  std_logic_vector(11 downto 0);
   -- timing of Y0: (c0, 0.550000ns)
signal Y1 :  std_logic_vector(11 downto 0);
   -- timing of Y1: (c0, 0.550000ns)
begin
   with X  select  Y0 <= 
      "000000001000" when "00000",
      "000001100100" when "00001",
      "000011000001" when "00010",
      "000100011101" when "00011",
      "000101111001" when "00100",
      "000111010110" when "00101",
      "001000110010" when "00110",
      "001010001110" when "00111",
      "001011101011" when "01000",
      "001101000111" when "01001",
      "001110100011" when "01010",
      "010000000000" when "01011",
      "010001011100" when "01100",
      "010010111000" when "01101",
      "010100010101" when "01110",
      "010101110001" when "01111",
      "010111001101" when "10000",
      "011000101010" when "10001",
      "011010000110" when "10010",
      "011011100010" when "10011",
      "011100111111" when "10100",
      "011110011011" when "10101",
      "011111110111" when "10110",
      "100001010100" when "10111",
      "100010110000" when "11000",
      "100100001100" when "11001",
      "100101101001" when "11010",
      "100111000101" when "11011",
      "101000100001" when "11100",
      "101001111110" when "11101",
      "101011011010" when "11110",
      "101100110110" when "11111",
      "------------" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                 FixRealKCM_Freq500_uid77_T1_Freq500_uid83
-- VHDL generated for DummyFPGA @ 500MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 2
-- Target frequency (MHz): 500
-- Input signals: X
-- Output signals: Y
--  approx. input signal timings: X: (c0, 0.000000ns)
--  approx. output signal timings: Y: (c0, 0.550000ns)

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity FixRealKCM_Freq500_uid77_T1_Freq500_uid83 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(6 downto 0)   );
end entity;

architecture arch of FixRealKCM_Freq500_uid77_T1_Freq500_uid83 is
signal Y0 :  std_logic_vector(6 downto 0);
   -- timing of Y0: (c0, 0.550000ns)
signal Y1 :  std_logic_vector(6 downto 0);
   -- timing of Y1: (c0, 0.550000ns)
begin
   with X  select  Y0 <= 
      "0000000" when "00000",
      "0000011" when "00001",
      "0000110" when "00010",
      "0001001" when "00011",
      "0001100" when "00100",
      "0001110" when "00101",
      "0010001" when "00110",
      "0010100" when "00111",
      "0010111" when "01000",
      "0011010" when "01001",
      "0011101" when "01010",
      "0100000" when "01011",
      "0100011" when "01100",
      "0100110" when "01101",
      "0101000" when "01110",
      "0101011" when "01111",
      "0101110" when "10000",
      "0110001" when "10001",
      "0110100" when "10010",
      "0110111" when "10011",
      "0111010" when "10100",
      "0111101" when "10101",
      "0111111" when "10110",
      "1000010" when "10111",
      "1000101" when "11000",
      "1001000" when "11001",
      "1001011" when "11010",
      "1001110" when "11011",
      "1010001" when "11100",
      "1010100" when "11101",
      "1010111" when "11110",
      "1011001" when "11111",
      "-------" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                 FixRealKCM_Freq500_uid89_T0_Freq500_uid92
-- VHDL generated for DummyFPGA @ 500MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 2
-- Target frequency (MHz): 500
-- Input signals: X
-- Output signals: Y
--  approx. input signal timings: X: (c0, 0.000000ns)
--  approx. output signal timings: Y: (c0, 0.550000ns)

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity FixRealKCM_Freq500_uid89_T0_Freq500_uid92 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(20 downto 0)   );
end entity;

architecture arch of FixRealKCM_Freq500_uid89_T0_Freq500_uid92 is
signal Y0 :  std_logic_vector(20 downto 0);
   -- timing of Y0: (c0, 0.550000ns)
signal Y1 :  std_logic_vector(20 downto 0);
   -- timing of Y1: (c0, 0.550000ns)
begin
   with X  select  Y0 <= 
      "000000000000000000000" when "00000",
      "000001011000101110010" when "00001",
      "000010110001011100100" when "00010",
      "000100001010001010110" when "00011",
      "000101100010111001000" when "00100",
      "000110111011100111010" when "00101",
      "001000010100010101101" when "00110",
      "001001101101000011111" when "00111",
      "001011000101110010001" when "01000",
      "001100011110100000011" when "01001",
      "001101110111001110101" when "01010",
      "001111001111111100111" when "01011",
      "010000101000101011001" when "01100",
      "010010000001011001011" when "01101",
      "010011011010000111101" when "01110",
      "010100110010110101111" when "01111",
      "010110001011100100001" when "10000",
      "010111100100010010100" when "10001",
      "011000111101000000110" when "10010",
      "011010010101101111000" when "10011",
      "011011101110011101010" when "10100",
      "011101000111001011100" when "10101",
      "011110011111111001110" when "10110",
      "011111111000101000000" when "10111",
      "100001010001010110010" when "11000",
      "100010101010000100100" when "11001",
      "100100000010110010110" when "11010",
      "100101011011100001001" when "11011",
      "100110110100001111011" when "11100",
      "101000001100111101101" when "11101",
      "101001100101101011111" when "11110",
      "101010111110011010001" when "11111",
      "---------------------" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                 FixRealKCM_Freq500_uid89_T1_Freq500_uid95
-- VHDL generated for DummyFPGA @ 500MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 2
-- Target frequency (MHz): 500
-- Input signals: X
-- Output signals: Y
--  approx. input signal timings: X: (c0, 0.000000ns)
--  approx. output signal timings: Y: (c0, 0.550000ns)

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity FixRealKCM_Freq500_uid89_T1_Freq500_uid95 is
    port (X : in  std_logic_vector(2 downto 0);
          Y : out  std_logic_vector(15 downto 0)   );
end entity;

architecture arch of FixRealKCM_Freq500_uid89_T1_Freq500_uid95 is
signal Y0 :  std_logic_vector(15 downto 0);
   -- timing of Y0: (c0, 0.550000ns)
signal Y1 :  std_logic_vector(15 downto 0);
   -- timing of Y1: (c0, 0.550000ns)
begin
   with X  select  Y0 <= 
      "0000000000000000" when "000",
      "0001011000101110" when "001",
      "0010110001011101" when "010",
      "0100001010001011" when "011",
      "0101100010111001" when "100",
      "0110111011100111" when "101",
      "1000010100010110" when "110",
      "1001101101000100" when "111",
      "----------------" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                     FixFunctionByTable_Freq500_uid104
-- Evaluator for exp(x*1b-1) on [-1,1) for lsbIn=-9 (wIn=10), msbout=0, lsbOut=-13 (wOut=14). Out interval: [0.606531; 1.64711]. Output is unsigned

-- VHDL generated for DummyFPGA @ 500MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin (2010-2018)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 2
-- Target frequency (MHz): 500
-- Input signals: X
-- Output signals: Y
--  approx. input signal timings: X: (c0, 0.000000ns)
--  approx. output signal timings: Y: (c0, 0.550000ns)

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity FixFunctionByTable_Freq500_uid104 is
    port (X : in  std_logic_vector(9 downto 0);
          Y : out  std_logic_vector(13 downto 0)   );
end entity;

architecture arch of FixFunctionByTable_Freq500_uid104 is
signal Y0 :  std_logic_vector(13 downto 0);
   -- timing of Y0: (c0, 0.550000ns)
signal Y1 :  std_logic_vector(13 downto 0);
   -- timing of Y1: (c0, 0.550000ns)
begin
   with X  select  Y0 <= 
      "10000000000000" when "0000000000",
      "10000000001000" when "0000000001",
      "10000000010000" when "0000000010",
      "10000000011000" when "0000000011",
      "10000000100000" when "0000000100",
      "10000000101000" when "0000000101",
      "10000000110000" when "0000000110",
      "10000000111000" when "0000000111",
      "10000001000000" when "0000001000",
      "10000001001000" when "0000001001",
      "10000001010000" when "0000001010",
      "10000001011000" when "0000001011",
      "10000001100001" when "0000001100",
      "10000001101001" when "0000001101",
      "10000001110001" when "0000001110",
      "10000001111001" when "0000001111",
      "10000010000001" when "0000010000",
      "10000010001001" when "0000010001",
      "10000010010001" when "0000010010",
      "10000010011001" when "0000010011",
      "10000010100010" when "0000010100",
      "10000010101010" when "0000010101",
      "10000010110010" when "0000010110",
      "10000010111010" when "0000010111",
      "10000011000010" when "0000011000",
      "10000011001010" when "0000011001",
      "10000011010011" when "0000011010",
      "10000011011011" when "0000011011",
      "10000011100011" when "0000011100",
      "10000011101011" when "0000011101",
      "10000011110100" when "0000011110",
      "10000011111100" when "0000011111",
      "10000100000100" when "0000100000",
      "10000100001100" when "0000100001",
      "10000100010101" when "0000100010",
      "10000100011101" when "0000100011",
      "10000100100101" when "0000100100",
      "10000100101101" when "0000100101",
      "10000100110110" when "0000100110",
      "10000100111110" when "0000100111",
      "10000101000110" when "0000101000",
      "10000101001111" when "0000101001",
      "10000101010111" when "0000101010",
      "10000101011111" when "0000101011",
      "10000101101000" when "0000101100",
      "10000101110000" when "0000101101",
      "10000101111000" when "0000101110",
      "10000110000001" when "0000101111",
      "10000110001001" when "0000110000",
      "10000110010010" when "0000110001",
      "10000110011010" when "0000110010",
      "10000110100010" when "0000110011",
      "10000110101011" when "0000110100",
      "10000110110011" when "0000110101",
      "10000110111100" when "0000110110",
      "10000111000100" when "0000110111",
      "10000111001100" when "0000111000",
      "10000111010101" when "0000111001",
      "10000111011101" when "0000111010",
      "10000111100110" when "0000111011",
      "10000111101110" when "0000111100",
      "10000111110111" when "0000111101",
      "10000111111111" when "0000111110",
      "10001000001000" when "0000111111",
      "10001000010000" when "0001000000",
      "10001000011001" when "0001000001",
      "10001000100001" when "0001000010",
      "10001000101010" when "0001000011",
      "10001000110010" when "0001000100",
      "10001000111011" when "0001000101",
      "10001001000100" when "0001000110",
      "10001001001100" when "0001000111",
      "10001001010101" when "0001001000",
      "10001001011101" when "0001001001",
      "10001001100110" when "0001001010",
      "10001001101111" when "0001001011",
      "10001001110111" when "0001001100",
      "10001010000000" when "0001001101",
      "10001010001000" when "0001001110",
      "10001010010001" when "0001001111",
      "10001010011010" when "0001010000",
      "10001010100010" when "0001010001",
      "10001010101011" when "0001010010",
      "10001010110100" when "0001010011",
      "10001010111100" when "0001010100",
      "10001011000101" when "0001010101",
      "10001011001110" when "0001010110",
      "10001011010110" when "0001010111",
      "10001011011111" when "0001011000",
      "10001011101000" when "0001011001",
      "10001011110001" when "0001011010",
      "10001011111001" when "0001011011",
      "10001100000010" when "0001011100",
      "10001100001011" when "0001011101",
      "10001100010100" when "0001011110",
      "10001100011100" when "0001011111",
      "10001100100101" when "0001100000",
      "10001100101110" when "0001100001",
      "10001100110111" when "0001100010",
      "10001101000000" when "0001100011",
      "10001101001000" when "0001100100",
      "10001101010001" when "0001100101",
      "10001101011010" when "0001100110",
      "10001101100011" when "0001100111",
      "10001101101100" when "0001101000",
      "10001101110101" when "0001101001",
      "10001101111101" when "0001101010",
      "10001110000110" when "0001101011",
      "10001110001111" when "0001101100",
      "10001110011000" when "0001101101",
      "10001110100001" when "0001101110",
      "10001110101010" when "0001101111",
      "10001110110011" when "0001110000",
      "10001110111100" when "0001110001",
      "10001111000101" when "0001110010",
      "10001111001110" when "0001110011",
      "10001111010111" when "0001110100",
      "10001111100000" when "0001110101",
      "10001111101001" when "0001110110",
      "10001111110010" when "0001110111",
      "10001111111011" when "0001111000",
      "10010000000100" when "0001111001",
      "10010000001101" when "0001111010",
      "10010000010110" when "0001111011",
      "10010000011111" when "0001111100",
      "10010000101000" when "0001111101",
      "10010000110001" when "0001111110",
      "10010000111010" when "0001111111",
      "10010001000011" when "0010000000",
      "10010001001100" when "0010000001",
      "10010001010101" when "0010000010",
      "10010001011110" when "0010000011",
      "10010001100111" when "0010000100",
      "10010001110000" when "0010000101",
      "10010001111001" when "0010000110",
      "10010010000010" when "0010000111",
      "10010010001100" when "0010001000",
      "10010010010101" when "0010001001",
      "10010010011110" when "0010001010",
      "10010010100111" when "0010001011",
      "10010010110000" when "0010001100",
      "10010010111001" when "0010001101",
      "10010011000011" when "0010001110",
      "10010011001100" when "0010001111",
      "10010011010101" when "0010010000",
      "10010011011110" when "0010010001",
      "10010011100111" when "0010010010",
      "10010011110001" when "0010010011",
      "10010011111010" when "0010010100",
      "10010100000011" when "0010010101",
      "10010100001100" when "0010010110",
      "10010100010110" when "0010010111",
      "10010100011111" when "0010011000",
      "10010100101000" when "0010011001",
      "10010100110001" when "0010011010",
      "10010100111011" when "0010011011",
      "10010101000100" when "0010011100",
      "10010101001101" when "0010011101",
      "10010101010111" when "0010011110",
      "10010101100000" when "0010011111",
      "10010101101001" when "0010100000",
      "10010101110011" when "0010100001",
      "10010101111100" when "0010100010",
      "10010110000110" when "0010100011",
      "10010110001111" when "0010100100",
      "10010110011000" when "0010100101",
      "10010110100010" when "0010100110",
      "10010110101011" when "0010100111",
      "10010110110101" when "0010101000",
      "10010110111110" when "0010101001",
      "10010111000111" when "0010101010",
      "10010111010001" when "0010101011",
      "10010111011010" when "0010101100",
      "10010111100100" when "0010101101",
      "10010111101101" when "0010101110",
      "10010111110111" when "0010101111",
      "10011000000000" when "0010110000",
      "10011000001010" when "0010110001",
      "10011000010011" when "0010110010",
      "10011000011101" when "0010110011",
      "10011000100110" when "0010110100",
      "10011000110000" when "0010110101",
      "10011000111001" when "0010110110",
      "10011001000011" when "0010110111",
      "10011001001101" when "0010111000",
      "10011001010110" when "0010111001",
      "10011001100000" when "0010111010",
      "10011001101001" when "0010111011",
      "10011001110011" when "0010111100",
      "10011001111101" when "0010111101",
      "10011010000110" when "0010111110",
      "10011010010000" when "0010111111",
      "10011010011001" when "0011000000",
      "10011010100011" when "0011000001",
      "10011010101101" when "0011000010",
      "10011010110110" when "0011000011",
      "10011011000000" when "0011000100",
      "10011011001010" when "0011000101",
      "10011011010100" when "0011000110",
      "10011011011101" when "0011000111",
      "10011011100111" when "0011001000",
      "10011011110001" when "0011001001",
      "10011011111010" when "0011001010",
      "10011100000100" when "0011001011",
      "10011100001110" when "0011001100",
      "10011100011000" when "0011001101",
      "10011100100001" when "0011001110",
      "10011100101011" when "0011001111",
      "10011100110101" when "0011010000",
      "10011100111111" when "0011010001",
      "10011101001001" when "0011010010",
      "10011101010010" when "0011010011",
      "10011101011100" when "0011010100",
      "10011101100110" when "0011010101",
      "10011101110000" when "0011010110",
      "10011101111010" when "0011010111",
      "10011110000100" when "0011011000",
      "10011110001110" when "0011011001",
      "10011110011000" when "0011011010",
      "10011110100001" when "0011011011",
      "10011110101011" when "0011011100",
      "10011110110101" when "0011011101",
      "10011110111111" when "0011011110",
      "10011111001001" when "0011011111",
      "10011111010011" when "0011100000",
      "10011111011101" when "0011100001",
      "10011111100111" when "0011100010",
      "10011111110001" when "0011100011",
      "10011111111011" when "0011100100",
      "10100000000101" when "0011100101",
      "10100000001111" when "0011100110",
      "10100000011001" when "0011100111",
      "10100000100011" when "0011101000",
      "10100000101101" when "0011101001",
      "10100000110111" when "0011101010",
      "10100001000001" when "0011101011",
      "10100001001011" when "0011101100",
      "10100001010101" when "0011101101",
      "10100001011111" when "0011101110",
      "10100001101010" when "0011101111",
      "10100001110100" when "0011110000",
      "10100001111110" when "0011110001",
      "10100010001000" when "0011110010",
      "10100010010010" when "0011110011",
      "10100010011100" when "0011110100",
      "10100010100110" when "0011110101",
      "10100010110001" when "0011110110",
      "10100010111011" when "0011110111",
      "10100011000101" when "0011111000",
      "10100011001111" when "0011111001",
      "10100011011001" when "0011111010",
      "10100011100100" when "0011111011",
      "10100011101110" when "0011111100",
      "10100011111000" when "0011111101",
      "10100100000010" when "0011111110",
      "10100100001100" when "0011111111",
      "10100100010111" when "0100000000",
      "10100100100001" when "0100000001",
      "10100100101011" when "0100000010",
      "10100100110110" when "0100000011",
      "10100101000000" when "0100000100",
      "10100101001010" when "0100000101",
      "10100101010101" when "0100000110",
      "10100101011111" when "0100000111",
      "10100101101001" when "0100001000",
      "10100101110100" when "0100001001",
      "10100101111110" when "0100001010",
      "10100110001000" when "0100001011",
      "10100110010011" when "0100001100",
      "10100110011101" when "0100001101",
      "10100110101000" when "0100001110",
      "10100110110010" when "0100001111",
      "10100110111100" when "0100010000",
      "10100111000111" when "0100010001",
      "10100111010001" when "0100010010",
      "10100111011100" when "0100010011",
      "10100111100110" when "0100010100",
      "10100111110001" when "0100010101",
      "10100111111011" when "0100010110",
      "10101000000110" when "0100010111",
      "10101000010000" when "0100011000",
      "10101000011011" when "0100011001",
      "10101000100101" when "0100011010",
      "10101000110000" when "0100011011",
      "10101000111010" when "0100011100",
      "10101001000101" when "0100011101",
      "10101001001111" when "0100011110",
      "10101001011010" when "0100011111",
      "10101001100101" when "0100100000",
      "10101001101111" when "0100100001",
      "10101001111010" when "0100100010",
      "10101010000100" when "0100100011",
      "10101010001111" when "0100100100",
      "10101010011010" when "0100100101",
      "10101010100100" when "0100100110",
      "10101010101111" when "0100100111",
      "10101010111010" when "0100101000",
      "10101011000100" when "0100101001",
      "10101011001111" when "0100101010",
      "10101011011010" when "0100101011",
      "10101011100101" when "0100101100",
      "10101011101111" when "0100101101",
      "10101011111010" when "0100101110",
      "10101100000101" when "0100101111",
      "10101100010000" when "0100110000",
      "10101100011010" when "0100110001",
      "10101100100101" when "0100110010",
      "10101100110000" when "0100110011",
      "10101100111011" when "0100110100",
      "10101101000101" when "0100110101",
      "10101101010000" when "0100110110",
      "10101101011011" when "0100110111",
      "10101101100110" when "0100111000",
      "10101101110001" when "0100111001",
      "10101101111100" when "0100111010",
      "10101110000111" when "0100111011",
      "10101110010001" when "0100111100",
      "10101110011100" when "0100111101",
      "10101110100111" when "0100111110",
      "10101110110010" when "0100111111",
      "10101110111101" when "0101000000",
      "10101111001000" when "0101000001",
      "10101111010011" when "0101000010",
      "10101111011110" when "0101000011",
      "10101111101001" when "0101000100",
      "10101111110100" when "0101000101",
      "10101111111111" when "0101000110",
      "10110000001010" when "0101000111",
      "10110000010101" when "0101001000",
      "10110000100000" when "0101001001",
      "10110000101011" when "0101001010",
      "10110000110110" when "0101001011",
      "10110001000001" when "0101001100",
      "10110001001100" when "0101001101",
      "10110001010111" when "0101001110",
      "10110001100010" when "0101001111",
      "10110001101101" when "0101010000",
      "10110001111001" when "0101010001",
      "10110010000100" when "0101010010",
      "10110010001111" when "0101010011",
      "10110010011010" when "0101010100",
      "10110010100101" when "0101010101",
      "10110010110000" when "0101010110",
      "10110010111011" when "0101010111",
      "10110011000111" when "0101011000",
      "10110011010010" when "0101011001",
      "10110011011101" when "0101011010",
      "10110011101000" when "0101011011",
      "10110011110100" when "0101011100",
      "10110011111111" when "0101011101",
      "10110100001010" when "0101011110",
      "10110100010101" when "0101011111",
      "10110100100001" when "0101100000",
      "10110100101100" when "0101100001",
      "10110100110111" when "0101100010",
      "10110101000010" when "0101100011",
      "10110101001110" when "0101100100",
      "10110101011001" when "0101100101",
      "10110101100100" when "0101100110",
      "10110101110000" when "0101100111",
      "10110101111011" when "0101101000",
      "10110110000111" when "0101101001",
      "10110110010010" when "0101101010",
      "10110110011101" when "0101101011",
      "10110110101001" when "0101101100",
      "10110110110100" when "0101101101",
      "10110111000000" when "0101101110",
      "10110111001011" when "0101101111",
      "10110111010110" when "0101110000",
      "10110111100010" when "0101110001",
      "10110111101101" when "0101110010",
      "10110111111001" when "0101110011",
      "10111000000100" when "0101110100",
      "10111000010000" when "0101110101",
      "10111000011011" when "0101110110",
      "10111000100111" when "0101110111",
      "10111000110011" when "0101111000",
      "10111000111110" when "0101111001",
      "10111001001010" when "0101111010",
      "10111001010101" when "0101111011",
      "10111001100001" when "0101111100",
      "10111001101100" when "0101111101",
      "10111001111000" when "0101111110",
      "10111010000100" when "0101111111",
      "10111010001111" when "0110000000",
      "10111010011011" when "0110000001",
      "10111010100111" when "0110000010",
      "10111010110010" when "0110000011",
      "10111010111110" when "0110000100",
      "10111011001010" when "0110000101",
      "10111011010101" when "0110000110",
      "10111011100001" when "0110000111",
      "10111011101101" when "0110001000",
      "10111011111001" when "0110001001",
      "10111100000100" when "0110001010",
      "10111100010000" when "0110001011",
      "10111100011100" when "0110001100",
      "10111100101000" when "0110001101",
      "10111100110011" when "0110001110",
      "10111100111111" when "0110001111",
      "10111101001011" when "0110010000",
      "10111101010111" when "0110010001",
      "10111101100011" when "0110010010",
      "10111101101111" when "0110010011",
      "10111101111010" when "0110010100",
      "10111110000110" when "0110010101",
      "10111110010010" when "0110010110",
      "10111110011110" when "0110010111",
      "10111110101010" when "0110011000",
      "10111110110110" when "0110011001",
      "10111111000010" when "0110011010",
      "10111111001110" when "0110011011",
      "10111111011010" when "0110011100",
      "10111111100110" when "0110011101",
      "10111111110010" when "0110011110",
      "10111111111110" when "0110011111",
      "11000000001010" when "0110100000",
      "11000000010110" when "0110100001",
      "11000000100010" when "0110100010",
      "11000000101110" when "0110100011",
      "11000000111010" when "0110100100",
      "11000001000110" when "0110100101",
      "11000001010010" when "0110100110",
      "11000001011110" when "0110100111",
      "11000001101010" when "0110101000",
      "11000001110110" when "0110101001",
      "11000010000010" when "0110101010",
      "11000010001110" when "0110101011",
      "11000010011011" when "0110101100",
      "11000010100111" when "0110101101",
      "11000010110011" when "0110101110",
      "11000010111111" when "0110101111",
      "11000011001011" when "0110110000",
      "11000011011000" when "0110110001",
      "11000011100100" when "0110110010",
      "11000011110000" when "0110110011",
      "11000011111100" when "0110110100",
      "11000100001000" when "0110110101",
      "11000100010101" when "0110110110",
      "11000100100001" when "0110110111",
      "11000100101101" when "0110111000",
      "11000100111010" when "0110111001",
      "11000101000110" when "0110111010",
      "11000101010010" when "0110111011",
      "11000101011111" when "0110111100",
      "11000101101011" when "0110111101",
      "11000101110111" when "0110111110",
      "11000110000100" when "0110111111",
      "11000110010000" when "0111000000",
      "11000110011100" when "0111000001",
      "11000110101001" when "0111000010",
      "11000110110101" when "0111000011",
      "11000111000010" when "0111000100",
      "11000111001110" when "0111000101",
      "11000111011011" when "0111000110",
      "11000111100111" when "0111000111",
      "11000111110100" when "0111001000",
      "11001000000000" when "0111001001",
      "11001000001101" when "0111001010",
      "11001000011001" when "0111001011",
      "11001000100110" when "0111001100",
      "11001000110010" when "0111001101",
      "11001000111111" when "0111001110",
      "11001001001011" when "0111001111",
      "11001001011000" when "0111010000",
      "11001001100100" when "0111010001",
      "11001001110001" when "0111010010",
      "11001001111110" when "0111010011",
      "11001010001010" when "0111010100",
      "11001010010111" when "0111010101",
      "11001010100100" when "0111010110",
      "11001010110000" when "0111010111",
      "11001010111101" when "0111011000",
      "11001011001010" when "0111011001",
      "11001011010110" when "0111011010",
      "11001011100011" when "0111011011",
      "11001011110000" when "0111011100",
      "11001011111100" when "0111011101",
      "11001100001001" when "0111011110",
      "11001100010110" when "0111011111",
      "11001100100011" when "0111100000",
      "11001100110000" when "0111100001",
      "11001100111100" when "0111100010",
      "11001101001001" when "0111100011",
      "11001101010110" when "0111100100",
      "11001101100011" when "0111100101",
      "11001101110000" when "0111100110",
      "11001101111101" when "0111100111",
      "11001110001001" when "0111101000",
      "11001110010110" when "0111101001",
      "11001110100011" when "0111101010",
      "11001110110000" when "0111101011",
      "11001110111101" when "0111101100",
      "11001111001010" when "0111101101",
      "11001111010111" when "0111101110",
      "11001111100100" when "0111101111",
      "11001111110001" when "0111110000",
      "11001111111110" when "0111110001",
      "11010000001011" when "0111110010",
      "11010000011000" when "0111110011",
      "11010000100101" when "0111110100",
      "11010000110010" when "0111110101",
      "11010000111111" when "0111110110",
      "11010001001100" when "0111110111",
      "11010001011001" when "0111111000",
      "11010001100110" when "0111111001",
      "11010001110011" when "0111111010",
      "11010010000001" when "0111111011",
      "11010010001110" when "0111111100",
      "11010010011011" when "0111111101",
      "11010010101000" when "0111111110",
      "11010010110101" when "0111111111",
      "01001101101001" when "1000000000",
      "01001101101110" when "1000000001",
      "01001101110010" when "1000000010",
      "01001101110111" when "1000000011",
      "01001101111100" when "1000000100",
      "01001110000001" when "1000000101",
      "01001110000110" when "1000000110",
      "01001110001011" when "1000000111",
      "01001110010000" when "1000001000",
      "01001110010101" when "1000001001",
      "01001110011001" when "1000001010",
      "01001110011110" when "1000001011",
      "01001110100011" when "1000001100",
      "01001110101000" when "1000001101",
      "01001110101101" when "1000001110",
      "01001110110010" when "1000001111",
      "01001110110111" when "1000010000",
      "01001110111100" when "1000010001",
      "01001111000001" when "1000010010",
      "01001111000110" when "1000010011",
      "01001111001011" when "1000010100",
      "01001111010000" when "1000010101",
      "01001111010101" when "1000010110",
      "01001111011010" when "1000010111",
      "01001111011111" when "1000011000",
      "01001111100011" when "1000011001",
      "01001111101000" when "1000011010",
      "01001111101101" when "1000011011",
      "01001111110010" when "1000011100",
      "01001111110111" when "1000011101",
      "01001111111100" when "1000011110",
      "01010000000001" when "1000011111",
      "01010000000110" when "1000100000",
      "01010000001011" when "1000100001",
      "01010000010000" when "1000100010",
      "01010000010101" when "1000100011",
      "01010000011010" when "1000100100",
      "01010000100000" when "1000100101",
      "01010000100101" when "1000100110",
      "01010000101010" when "1000100111",
      "01010000101111" when "1000101000",
      "01010000110100" when "1000101001",
      "01010000111001" when "1000101010",
      "01010000111110" when "1000101011",
      "01010001000011" when "1000101100",
      "01010001001000" when "1000101101",
      "01010001001101" when "1000101110",
      "01010001010010" when "1000101111",
      "01010001010111" when "1000110000",
      "01010001011100" when "1000110001",
      "01010001100001" when "1000110010",
      "01010001100110" when "1000110011",
      "01010001101100" when "1000110100",
      "01010001110001" when "1000110101",
      "01010001110110" when "1000110110",
      "01010001111011" when "1000110111",
      "01010010000000" when "1000111000",
      "01010010000101" when "1000111001",
      "01010010001010" when "1000111010",
      "01010010001111" when "1000111011",
      "01010010010101" when "1000111100",
      "01010010011010" when "1000111101",
      "01010010011111" when "1000111110",
      "01010010100100" when "1000111111",
      "01010010101001" when "1001000000",
      "01010010101110" when "1001000001",
      "01010010110011" when "1001000010",
      "01010010111001" when "1001000011",
      "01010010111110" when "1001000100",
      "01010011000011" when "1001000101",
      "01010011001000" when "1001000110",
      "01010011001101" when "1001000111",
      "01010011010011" when "1001001000",
      "01010011011000" when "1001001001",
      "01010011011101" when "1001001010",
      "01010011100010" when "1001001011",
      "01010011100111" when "1001001100",
      "01010011101101" when "1001001101",
      "01010011110010" when "1001001110",
      "01010011110111" when "1001001111",
      "01010011111100" when "1001010000",
      "01010100000010" when "1001010001",
      "01010100000111" when "1001010010",
      "01010100001100" when "1001010011",
      "01010100010001" when "1001010100",
      "01010100010111" when "1001010101",
      "01010100011100" when "1001010110",
      "01010100100001" when "1001010111",
      "01010100100111" when "1001011000",
      "01010100101100" when "1001011001",
      "01010100110001" when "1001011010",
      "01010100110110" when "1001011011",
      "01010100111100" when "1001011100",
      "01010101000001" when "1001011101",
      "01010101000110" when "1001011110",
      "01010101001100" when "1001011111",
      "01010101010001" when "1001100000",
      "01010101010110" when "1001100001",
      "01010101011100" when "1001100010",
      "01010101100001" when "1001100011",
      "01010101100110" when "1001100100",
      "01010101101100" when "1001100101",
      "01010101110001" when "1001100110",
      "01010101110110" when "1001100111",
      "01010101111100" when "1001101000",
      "01010110000001" when "1001101001",
      "01010110000111" when "1001101010",
      "01010110001100" when "1001101011",
      "01010110010001" when "1001101100",
      "01010110010111" when "1001101101",
      "01010110011100" when "1001101110",
      "01010110100010" when "1001101111",
      "01010110100111" when "1001110000",
      "01010110101100" when "1001110001",
      "01010110110010" when "1001110010",
      "01010110110111" when "1001110011",
      "01010110111101" when "1001110100",
      "01010111000010" when "1001110101",
      "01010111001000" when "1001110110",
      "01010111001101" when "1001110111",
      "01010111010010" when "1001111000",
      "01010111011000" when "1001111001",
      "01010111011101" when "1001111010",
      "01010111100011" when "1001111011",
      "01010111101000" when "1001111100",
      "01010111101110" when "1001111101",
      "01010111110011" when "1001111110",
      "01010111111001" when "1001111111",
      "01010111111110" when "1010000000",
      "01011000000100" when "1010000001",
      "01011000001001" when "1010000010",
      "01011000001111" when "1010000011",
      "01011000010100" when "1010000100",
      "01011000011010" when "1010000101",
      "01011000011111" when "1010000110",
      "01011000100101" when "1010000111",
      "01011000101010" when "1010001000",
      "01011000110000" when "1010001001",
      "01011000110110" when "1010001010",
      "01011000111011" when "1010001011",
      "01011001000001" when "1010001100",
      "01011001000110" when "1010001101",
      "01011001001100" when "1010001110",
      "01011001010001" when "1010001111",
      "01011001010111" when "1010010000",
      "01011001011101" when "1010010001",
      "01011001100010" when "1010010010",
      "01011001101000" when "1010010011",
      "01011001101101" when "1010010100",
      "01011001110011" when "1010010101",
      "01011001111001" when "1010010110",
      "01011001111110" when "1010010111",
      "01011010000100" when "1010011000",
      "01011010001001" when "1010011001",
      "01011010001111" when "1010011010",
      "01011010010101" when "1010011011",
      "01011010011010" when "1010011100",
      "01011010100000" when "1010011101",
      "01011010100110" when "1010011110",
      "01011010101011" when "1010011111",
      "01011010110001" when "1010100000",
      "01011010110111" when "1010100001",
      "01011010111100" when "1010100010",
      "01011011000010" when "1010100011",
      "01011011001000" when "1010100100",
      "01011011001101" when "1010100101",
      "01011011010011" when "1010100110",
      "01011011011001" when "1010100111",
      "01011011011111" when "1010101000",
      "01011011100100" when "1010101001",
      "01011011101010" when "1010101010",
      "01011011110000" when "1010101011",
      "01011011110101" when "1010101100",
      "01011011111011" when "1010101101",
      "01011100000001" when "1010101110",
      "01011100000111" when "1010101111",
      "01011100001100" when "1010110000",
      "01011100010010" when "1010110001",
      "01011100011000" when "1010110010",
      "01011100011110" when "1010110011",
      "01011100100100" when "1010110100",
      "01011100101001" when "1010110101",
      "01011100101111" when "1010110110",
      "01011100110101" when "1010110111",
      "01011100111011" when "1010111000",
      "01011101000001" when "1010111001",
      "01011101000110" when "1010111010",
      "01011101001100" when "1010111011",
      "01011101010010" when "1010111100",
      "01011101011000" when "1010111101",
      "01011101011110" when "1010111110",
      "01011101100100" when "1010111111",
      "01011101101001" when "1011000000",
      "01011101101111" when "1011000001",
      "01011101110101" when "1011000010",
      "01011101111011" when "1011000011",
      "01011110000001" when "1011000100",
      "01011110000111" when "1011000101",
      "01011110001101" when "1011000110",
      "01011110010011" when "1011000111",
      "01011110011000" when "1011001000",
      "01011110011110" when "1011001001",
      "01011110100100" when "1011001010",
      "01011110101010" when "1011001011",
      "01011110110000" when "1011001100",
      "01011110110110" when "1011001101",
      "01011110111100" when "1011001110",
      "01011111000010" when "1011001111",
      "01011111001000" when "1011010000",
      "01011111001110" when "1011010001",
      "01011111010100" when "1011010010",
      "01011111011010" when "1011010011",
      "01011111100000" when "1011010100",
      "01011111100110" when "1011010101",
      "01011111101100" when "1011010110",
      "01011111110010" when "1011010111",
      "01011111111000" when "1011011000",
      "01011111111110" when "1011011001",
      "01100000000100" when "1011011010",
      "01100000001010" when "1011011011",
      "01100000010000" when "1011011100",
      "01100000010110" when "1011011101",
      "01100000011100" when "1011011110",
      "01100000100010" when "1011011111",
      "01100000101000" when "1011100000",
      "01100000101110" when "1011100001",
      "01100000110100" when "1011100010",
      "01100000111010" when "1011100011",
      "01100001000000" when "1011100100",
      "01100001000110" when "1011100101",
      "01100001001100" when "1011100110",
      "01100001010010" when "1011100111",
      "01100001011000" when "1011101000",
      "01100001011110" when "1011101001",
      "01100001100100" when "1011101010",
      "01100001101010" when "1011101011",
      "01100001110001" when "1011101100",
      "01100001110111" when "1011101101",
      "01100001111101" when "1011101110",
      "01100010000011" when "1011101111",
      "01100010001001" when "1011110000",
      "01100010001111" when "1011110001",
      "01100010010101" when "1011110010",
      "01100010011011" when "1011110011",
      "01100010100010" when "1011110100",
      "01100010101000" when "1011110101",
      "01100010101110" when "1011110110",
      "01100010110100" when "1011110111",
      "01100010111010" when "1011111000",
      "01100011000000" when "1011111001",
      "01100011000111" when "1011111010",
      "01100011001101" when "1011111011",
      "01100011010011" when "1011111100",
      "01100011011001" when "1011111101",
      "01100011011111" when "1011111110",
      "01100011100110" when "1011111111",
      "01100011101100" when "1100000000",
      "01100011110010" when "1100000001",
      "01100011111000" when "1100000010",
      "01100011111111" when "1100000011",
      "01100100000101" when "1100000100",
      "01100100001011" when "1100000101",
      "01100100010001" when "1100000110",
      "01100100011000" when "1100000111",
      "01100100011110" when "1100001000",
      "01100100100100" when "1100001001",
      "01100100101011" when "1100001010",
      "01100100110001" when "1100001011",
      "01100100110111" when "1100001100",
      "01100100111101" when "1100001101",
      "01100101000100" when "1100001110",
      "01100101001010" when "1100001111",
      "01100101010000" when "1100010000",
      "01100101010111" when "1100010001",
      "01100101011101" when "1100010010",
      "01100101100011" when "1100010011",
      "01100101101010" when "1100010100",
      "01100101110000" when "1100010101",
      "01100101110110" when "1100010110",
      "01100101111101" when "1100010111",
      "01100110000011" when "1100011000",
      "01100110001010" when "1100011001",
      "01100110010000" when "1100011010",
      "01100110010110" when "1100011011",
      "01100110011101" when "1100011100",
      "01100110100011" when "1100011101",
      "01100110101010" when "1100011110",
      "01100110110000" when "1100011111",
      "01100110110110" when "1100100000",
      "01100110111101" when "1100100001",
      "01100111000011" when "1100100010",
      "01100111001010" when "1100100011",
      "01100111010000" when "1100100100",
      "01100111010111" when "1100100101",
      "01100111011101" when "1100100110",
      "01100111100100" when "1100100111",
      "01100111101010" when "1100101000",
      "01100111110001" when "1100101001",
      "01100111110111" when "1100101010",
      "01100111111110" when "1100101011",
      "01101000000100" when "1100101100",
      "01101000001011" when "1100101101",
      "01101000010001" when "1100101110",
      "01101000011000" when "1100101111",
      "01101000011110" when "1100110000",
      "01101000100101" when "1100110001",
      "01101000101011" when "1100110010",
      "01101000110010" when "1100110011",
      "01101000111000" when "1100110100",
      "01101000111111" when "1100110101",
      "01101001000101" when "1100110110",
      "01101001001100" when "1100110111",
      "01101001010011" when "1100111000",
      "01101001011001" when "1100111001",
      "01101001100000" when "1100111010",
      "01101001100110" when "1100111011",
      "01101001101101" when "1100111100",
      "01101001110100" when "1100111101",
      "01101001111010" when "1100111110",
      "01101010000001" when "1100111111",
      "01101010000111" when "1101000000",
      "01101010001110" when "1101000001",
      "01101010010101" when "1101000010",
      "01101010011011" when "1101000011",
      "01101010100010" when "1101000100",
      "01101010101001" when "1101000101",
      "01101010101111" when "1101000110",
      "01101010110110" when "1101000111",
      "01101010111101" when "1101001000",
      "01101011000011" when "1101001001",
      "01101011001010" when "1101001010",
      "01101011010001" when "1101001011",
      "01101011010111" when "1101001100",
      "01101011011110" when "1101001101",
      "01101011100101" when "1101001110",
      "01101011101100" when "1101001111",
      "01101011110010" when "1101010000",
      "01101011111001" when "1101010001",
      "01101100000000" when "1101010010",
      "01101100000111" when "1101010011",
      "01101100001101" when "1101010100",
      "01101100010100" when "1101010101",
      "01101100011011" when "1101010110",
      "01101100100010" when "1101010111",
      "01101100101000" when "1101011000",
      "01101100101111" when "1101011001",
      "01101100110110" when "1101011010",
      "01101100111101" when "1101011011",
      "01101101000100" when "1101011100",
      "01101101001010" when "1101011101",
      "01101101010001" when "1101011110",
      "01101101011000" when "1101011111",
      "01101101011111" when "1101100000",
      "01101101100110" when "1101100001",
      "01101101101101" when "1101100010",
      "01101101110100" when "1101100011",
      "01101101111010" when "1101100100",
      "01101110000001" when "1101100101",
      "01101110001000" when "1101100110",
      "01101110001111" when "1101100111",
      "01101110010110" when "1101101000",
      "01101110011101" when "1101101001",
      "01101110100100" when "1101101010",
      "01101110101011" when "1101101011",
      "01101110110010" when "1101101100",
      "01101110111001" when "1101101101",
      "01101110111111" when "1101101110",
      "01101111000110" when "1101101111",
      "01101111001101" when "1101110000",
      "01101111010100" when "1101110001",
      "01101111011011" when "1101110010",
      "01101111100010" when "1101110011",
      "01101111101001" when "1101110100",
      "01101111110000" when "1101110101",
      "01101111110111" when "1101110110",
      "01101111111110" when "1101110111",
      "01110000000101" when "1101111000",
      "01110000001100" when "1101111001",
      "01110000010011" when "1101111010",
      "01110000011010" when "1101111011",
      "01110000100001" when "1101111100",
      "01110000101000" when "1101111101",
      "01110000101111" when "1101111110",
      "01110000110110" when "1101111111",
      "01110000111101" when "1110000000",
      "01110001000100" when "1110000001",
      "01110001001100" when "1110000010",
      "01110001010011" when "1110000011",
      "01110001011010" when "1110000100",
      "01110001100001" when "1110000101",
      "01110001101000" when "1110000110",
      "01110001101111" when "1110000111",
      "01110001110110" when "1110001000",
      "01110001111101" when "1110001001",
      "01110010000100" when "1110001010",
      "01110010001011" when "1110001011",
      "01110010010011" when "1110001100",
      "01110010011010" when "1110001101",
      "01110010100001" when "1110001110",
      "01110010101000" when "1110001111",
      "01110010101111" when "1110010000",
      "01110010110110" when "1110010001",
      "01110010111110" when "1110010010",
      "01110011000101" when "1110010011",
      "01110011001100" when "1110010100",
      "01110011010011" when "1110010101",
      "01110011011010" when "1110010110",
      "01110011100010" when "1110010111",
      "01110011101001" when "1110011000",
      "01110011110000" when "1110011001",
      "01110011110111" when "1110011010",
      "01110011111111" when "1110011011",
      "01110100000110" when "1110011100",
      "01110100001101" when "1110011101",
      "01110100010100" when "1110011110",
      "01110100011100" when "1110011111",
      "01110100100011" when "1110100000",
      "01110100101010" when "1110100001",
      "01110100110001" when "1110100010",
      "01110100111001" when "1110100011",
      "01110101000000" when "1110100100",
      "01110101000111" when "1110100101",
      "01110101001111" when "1110100110",
      "01110101010110" when "1110100111",
      "01110101011101" when "1110101000",
      "01110101100101" when "1110101001",
      "01110101101100" when "1110101010",
      "01110101110011" when "1110101011",
      "01110101111011" when "1110101100",
      "01110110000010" when "1110101101",
      "01110110001010" when "1110101110",
      "01110110010001" when "1110101111",
      "01110110011000" when "1110110000",
      "01110110100000" when "1110110001",
      "01110110100111" when "1110110010",
      "01110110101111" when "1110110011",
      "01110110110110" when "1110110100",
      "01110110111101" when "1110110101",
      "01110111000101" when "1110110110",
      "01110111001100" when "1110110111",
      "01110111010100" when "1110111000",
      "01110111011011" when "1110111001",
      "01110111100011" when "1110111010",
      "01110111101010" when "1110111011",
      "01110111110010" when "1110111100",
      "01110111111001" when "1110111101",
      "01111000000001" when "1110111110",
      "01111000001000" when "1110111111",
      "01111000010000" when "1111000000",
      "01111000010111" when "1111000001",
      "01111000011111" when "1111000010",
      "01111000100110" when "1111000011",
      "01111000101110" when "1111000100",
      "01111000110101" when "1111000101",
      "01111000111101" when "1111000110",
      "01111001000100" when "1111000111",
      "01111001001100" when "1111001000",
      "01111001010100" when "1111001001",
      "01111001011011" when "1111001010",
      "01111001100011" when "1111001011",
      "01111001101010" when "1111001100",
      "01111001110010" when "1111001101",
      "01111001111010" when "1111001110",
      "01111010000001" when "1111001111",
      "01111010001001" when "1111010000",
      "01111010010000" when "1111010001",
      "01111010011000" when "1111010010",
      "01111010100000" when "1111010011",
      "01111010100111" when "1111010100",
      "01111010101111" when "1111010101",
      "01111010110111" when "1111010110",
      "01111010111110" when "1111010111",
      "01111011000110" when "1111011000",
      "01111011001110" when "1111011001",
      "01111011010110" when "1111011010",
      "01111011011101" when "1111011011",
      "01111011100101" when "1111011100",
      "01111011101101" when "1111011101",
      "01111011110100" when "1111011110",
      "01111011111100" when "1111011111",
      "01111100000100" when "1111100000",
      "01111100001100" when "1111100001",
      "01111100010011" when "1111100010",
      "01111100011011" when "1111100011",
      "01111100100011" when "1111100100",
      "01111100101011" when "1111100101",
      "01111100110011" when "1111100110",
      "01111100111010" when "1111100111",
      "01111101000010" when "1111101000",
      "01111101001010" when "1111101001",
      "01111101010010" when "1111101010",
      "01111101011010" when "1111101011",
      "01111101100010" when "1111101100",
      "01111101101001" when "1111101101",
      "01111101110001" when "1111101110",
      "01111101111001" when "1111101111",
      "01111110000001" when "1111110000",
      "01111110001001" when "1111110001",
      "01111110010001" when "1111110010",
      "01111110011001" when "1111110011",
      "01111110100001" when "1111110100",
      "01111110101000" when "1111110101",
      "01111110110000" when "1111110110",
      "01111110111000" when "1111110111",
      "01111111000000" when "1111111000",
      "01111111001000" when "1111111001",
      "01111111010000" when "1111111010",
      "01111111011000" when "1111111011",
      "01111111100000" when "1111111100",
      "01111111101000" when "1111111101",
      "01111111110000" when "1111111110",
      "01111111111000" when "1111111111",
      "--------------" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                     FixFunctionByTable_Freq500_uid107
-- Evaluator for (exp(x*1b-11)-1) on [-1,1) for lsbIn=-2 (wIn=3), msbout=-11, lsbOut=-13 (wOut=3). Out interval: [-0.000488162; 0.000366278]. Output is signed

-- VHDL generated for DummyFPGA @ 500MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin (2010-2018)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 2
-- Target frequency (MHz): 500
-- Input signals: X
-- Output signals: Y
--  approx. input signal timings: X: (c0, 0.000000ns)
--  approx. output signal timings: Y: (c0, 0.550000ns)

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity FixFunctionByTable_Freq500_uid107 is
    port (X : in  std_logic_vector(2 downto 0);
          Y : out  std_logic_vector(2 downto 0)   );
end entity;

architecture arch of FixFunctionByTable_Freq500_uid107 is
signal Y0 :  std_logic_vector(2 downto 0);
   -- timing of Y0: (c0, 0.550000ns)
signal Y1 :  std_logic_vector(2 downto 0);
   -- timing of Y1: (c0, 0.550000ns)
begin
   with X  select  Y0 <= 
      "000" when "000",
      "001" when "001",
      "010" when "010",
      "011" when "011",
      "100" when "100",
      "101" when "101",
      "110" when "110",
      "111" when "111",
      "---" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          IntAdder_19_Freq500_uid5
-- VHDL generated for DummyFPGA @ 500MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin (2008-2016)
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 2
-- Target frequency (MHz): 500
-- Input signals: X Y Cin
-- Output signals: R
--  approx. input signal timings: X: (c0, 0.000000ns)Y: (c0, 0.000000ns)Cin: (c0, 0.000000ns)
--  approx. output signal timings: R: (c0, 1.180000ns)

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntAdder_19_Freq500_uid5 is
    port (clk : in std_logic;
          X : in  std_logic_vector(18 downto 0);
          Y : in  std_logic_vector(18 downto 0);
          Cin : in  std_logic;
          R : out  std_logic_vector(18 downto 0)   );
end entity;

architecture arch of IntAdder_19_Freq500_uid5 is
signal Rtmp :  std_logic_vector(18 downto 0);
   -- timing of Rtmp: (c0, 1.180000ns)
begin
   Rtmp <= X + Y + Cin;
   R <= Rtmp;
end architecture;

--------------------------------------------------------------------------------
--                            LZC_10_Freq500_uid7
-- VHDL generated for DummyFPGA @ 500MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007)
--------------------------------------------------------------------------------
-- Pipeline depth: 1 cycles
-- Clock period (ns): 2
-- Target frequency (MHz): 500
-- Input signals: I
-- Output signals: O
--  approx. input signal timings: I: (c0, 0.000000ns)
--  approx. output signal timings: O: (c1, 0.980000ns)

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity LZC_10_Freq500_uid7 is
    port (clk : in std_logic;
          I : in  std_logic_vector(9 downto 0);
          O : out  std_logic_vector(3 downto 0)   );
end entity;

architecture arch of LZC_10_Freq500_uid7 is
signal level4 :  std_logic_vector(14 downto 0);
   -- timing of level4: (c0, 0.000000ns)
signal digit3 :  std_logic;
   -- timing of digit3: (c0, 0.570000ns)
signal level3, level3_d1 :  std_logic_vector(6 downto 0);
   -- timing of level3: (c0, 1.120000ns)
signal digit2, digit2_d1 :  std_logic;
   -- timing of digit2: (c0, 1.680000ns)
signal level2 :  std_logic_vector(2 downto 0);
   -- timing of level2: (c1, 0.430000ns)
signal lowBits :  std_logic_vector(1 downto 0);
   -- timing of lowBits: (c1, 0.980000ns)
signal outHighBits, outHighBits_d1 :  std_logic_vector(1 downto 0);
   -- timing of outHighBits: (c0, 1.680000ns)
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            level3_d1 <=  level3;
            digit2_d1 <=  digit2;
            outHighBits_d1 <=  outHighBits;
         end if;
      end process;
   -- pad input to the next power of two minus 1
   level4 <= I & "11111";
   -- Main iteration for large inputs
   digit3<= '1' when level4(14 downto 7) = "00000000" else '0';
   level3<= level4(6 downto 0) when digit3='1' else level4(14 downto 8);
   digit2<= '1' when level3(6 downto 3) = "0000" else '0';
   level2<= level3_d1(2 downto 0) when digit2_d1='1' else level3_d1(6 downto 4);
   -- Finish counting with one LUT
   with level2  select  lowBits <= 
      "11" when "000",
      "10" when "001",
      "01" when "010",
      "01" when "011",
      "00" when others;
   outHighBits <= digit3 & digit2 & "";
   O <= outHighBits_d1 & lowBits ;
end architecture;

--------------------------------------------------------------------------------
--                           LZOC_20_Freq500_uid11
-- VHDL generated for DummyFPGA @ 500MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007)
--------------------------------------------------------------------------------
-- Pipeline depth: 3 cycles
-- Clock period (ns): 2
-- Target frequency (MHz): 500
-- Input signals: I OZB
-- Output signals: O
--  approx. input signal timings: I: (c0, 0.550000ns)OZB: (c0, 0.000000ns)
--  approx. output signal timings: O: (c3, 0.410000ns)

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity LZOC_20_Freq500_uid11 is
    port (clk : in std_logic;
          I : in  std_logic_vector(19 downto 0);
          OZB : in  std_logic;
          O : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of LZOC_20_Freq500_uid11 is
signal sozb, sozb_d1, sozb_d2 :  std_logic;
   -- timing of sozb: (c0, 0.000000ns)
signal level5, level5_d1 :  std_logic_vector(30 downto 0);
   -- timing of level5: (c0, 0.550000ns)
signal digit4, digit4_d1, digit4_d2 :  std_logic;
   -- timing of digit4: (c0, 1.590000ns)
signal level4, level4_d1 :  std_logic_vector(14 downto 0);
   -- timing of level4: (c1, 0.340000ns)
signal digit3, digit3_d1 :  std_logic;
   -- timing of digit3: (c1, 1.360000ns)
signal level3 :  std_logic_vector(6 downto 0);
   -- timing of level3: (c2, 0.110000ns)
signal digit2 :  std_logic;
   -- timing of digit2: (c2, 1.110000ns)
signal level2, level2_d1 :  std_logic_vector(2 downto 0);
   -- timing of level2: (c2, 1.660000ns)
signal z :  std_logic_vector(2 downto 0);
   -- timing of z: (c3, 0.410000ns)
signal lowBits :  std_logic_vector(1 downto 0);
   -- timing of lowBits: (c3, 0.410000ns)
signal outHighBits, outHighBits_d1 :  std_logic_vector(2 downto 0);
   -- timing of outHighBits: (c2, 1.110000ns)
signal OZB_d1, OZB_d2, OZB_d3 :  std_logic;
   -- timing of OZB: (c0, 0.000000ns)
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            sozb_d1 <=  sozb;
            sozb_d2 <=  sozb_d1;
            level5_d1 <=  level5;
            digit4_d1 <=  digit4;
            digit4_d2 <=  digit4_d1;
            level4_d1 <=  level4;
            digit3_d1 <=  digit3;
            level2_d1 <=  level2;
            outHighBits_d1 <=  outHighBits;
            OZB_d1 <=  OZB;
            OZB_d2 <=  OZB_d1;
            OZB_d3 <=  OZB_d2;
         end if;
      end process;
   sozb <= OZB;
   -- pad input to the next power of two minus 1
   level5 <= I & (10 downto 0 => not sozb);
   -- Main iteration for large inputs
   digit4<= '1' when level5(30 downto 15) = (15 downto 0 => sozb) else '0';
   level4<= level5_d1(14 downto 0) when digit4_d1='1' else level5_d1(30 downto 16);
   digit3<= '1' when level4(14 downto 7) = (7 downto 0 => sozb_d1) else '0';
   level3<= level4_d1(6 downto 0) when digit3_d1='1' else level4_d1(14 downto 8);
   digit2<= '1' when level3(6 downto 3) = (3 downto 0 => sozb_d2) else '0';
   level2<= level3(2 downto 0) when digit2='1' else level3(6 downto 4);
   -- Finish counting with one LUT
   z <= level2_d1 when OZB_d3='0' else (not level2_d1);
   with z  select  lowBits <= 
      "11" when "000",
      "10" when "001",
      "01" when "010",
      "01" when "011",
      "00" when others;
   outHighBits <= digit4_d2 & digit3_d1 & digit2 & "";
   O <= outHighBits_d1 & lowBits ;
end architecture;

--------------------------------------------------------------------------------
--                   LeftShifter11_by_max_11_Freq500_uid13
-- VHDL generated for DummyFPGA @ 500MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca (2008-2011), Florent de Dinechin (2008-2019)
--------------------------------------------------------------------------------
-- Pipeline depth: 4 cycles
-- Clock period (ns): 2
-- Target frequency (MHz): 500
-- Input signals: X S
-- Output signals: R
--  approx. input signal timings: X: (c0, 1.650000ns)S: (c3, 1.460000ns)
--  approx. output signal timings: R: (c4, 1.375385ns)

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity LeftShifter11_by_max_11_Freq500_uid13 is
    port (clk : in std_logic;
          X : in  std_logic_vector(10 downto 0);
          S : in  std_logic_vector(3 downto 0);
          R : out  std_logic_vector(21 downto 0)   );
end entity;

architecture arch of LeftShifter11_by_max_11_Freq500_uid13 is
signal ps, ps_d1 :  std_logic_vector(3 downto 0);
   -- timing of ps: (c3, 1.460000ns)
signal level0, level0_d1, level0_d2, level0_d3 :  std_logic_vector(10 downto 0);
   -- timing of level0: (c0, 1.650000ns)
signal level1, level1_d1 :  std_logic_vector(11 downto 0);
   -- timing of level1: (c3, 1.460000ns)
signal level2 :  std_logic_vector(13 downto 0);
   -- timing of level2: (c4, 0.425385ns)
signal level3 :  std_logic_vector(17 downto 0);
   -- timing of level3: (c4, 0.425385ns)
signal level4 :  std_logic_vector(25 downto 0);
   -- timing of level4: (c4, 1.375385ns)
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            ps_d1 <=  ps;
            level0_d1 <=  level0;
            level0_d2 <=  level0_d1;
            level0_d3 <=  level0_d2;
            level1_d1 <=  level1;
         end if;
      end process;
   ps<= S;
   level0<= X;
   level1<= level0_d3 & (0 downto 0 => '0') when ps(0)= '1' else     (0 downto 0 => '0') & level0_d3;
   level2<= level1_d1 & (1 downto 0 => '0') when ps_d1(1)= '1' else     (1 downto 0 => '0') & level1_d1;
   level3<= level2 & (3 downto 0 => '0') when ps_d1(2)= '1' else     (3 downto 0 => '0') & level2;
   level4<= level3 & (7 downto 0 => '0') when ps_d1(3)= '1' else     (7 downto 0 => '0') & level3;
   R <= level4(21 downto 0);
end architecture;

--------------------------------------------------------------------------------
--                         IntAdder_24_Freq500_uid19
-- VHDL generated for DummyFPGA @ 500MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin (2008-2016)
--------------------------------------------------------------------------------
-- Pipeline depth: 2 cycles
-- Clock period (ns): 2
-- Target frequency (MHz): 500
-- Input signals: X Y Cin
-- Output signals: R
--  approx. input signal timings: X: (c1, 0.600000ns)Y: (c1, 1.150000ns)Cin: (c0, 0.000000ns)
--  approx. output signal timings: R: (c2, 0.590000ns)

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntAdder_24_Freq500_uid19 is
    port (clk : in std_logic;
          X : in  std_logic_vector(23 downto 0);
          Y : in  std_logic_vector(23 downto 0);
          Cin : in  std_logic;
          R : out  std_logic_vector(23 downto 0)   );
end entity;

architecture arch of IntAdder_24_Freq500_uid19 is
signal Cin_1, Cin_1_d1, Cin_1_d2 :  std_logic;
   -- timing of Cin_1: (c0, 0.000000ns)
signal X_1, X_1_d1 :  std_logic_vector(24 downto 0);
   -- timing of X_1: (c1, 0.600000ns)
signal Y_1, Y_1_d1 :  std_logic_vector(24 downto 0);
   -- timing of Y_1: (c1, 1.150000ns)
signal S_1 :  std_logic_vector(24 downto 0);
   -- timing of S_1: (c2, 0.590000ns)
signal R_1 :  std_logic_vector(23 downto 0);
   -- timing of R_1: (c2, 0.590000ns)
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            Cin_1_d1 <=  Cin_1;
            Cin_1_d2 <=  Cin_1_d1;
            X_1_d1 <=  X_1;
            Y_1_d1 <=  Y_1;
         end if;
      end process;
   Cin_1 <= Cin;
   X_1 <= '0' & X(23 downto 0);
   Y_1 <= '0' & Y(23 downto 0);
   S_1 <= X_1_d1 + Y_1_d1 + Cin_1_d2;
   R_1 <= S_1(23 downto 0);
   R <= R_1 ;
end architecture;

--------------------------------------------------------------------------------
--                         IntAdder_24_Freq500_uid22
-- VHDL generated for DummyFPGA @ 500MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin (2008-2016)
--------------------------------------------------------------------------------
-- Pipeline depth: 3 cycles
-- Clock period (ns): 2
-- Target frequency (MHz): 500
-- Input signals: X Y Cin
-- Output signals: R
--  approx. input signal timings: X: (c2, 0.590000ns)Y: (c2, 1.180000ns)Cin: (c0, 0.000000ns)
--  approx. output signal timings: R: (c3, 0.620000ns)

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntAdder_24_Freq500_uid22 is
    port (clk : in std_logic;
          X : in  std_logic_vector(23 downto 0);
          Y : in  std_logic_vector(23 downto 0);
          Cin : in  std_logic;
          R : out  std_logic_vector(23 downto 0)   );
end entity;

architecture arch of IntAdder_24_Freq500_uid22 is
signal Cin_1, Cin_1_d1, Cin_1_d2, Cin_1_d3 :  std_logic;
   -- timing of Cin_1: (c0, 0.000000ns)
signal X_1, X_1_d1 :  std_logic_vector(24 downto 0);
   -- timing of X_1: (c2, 0.590000ns)
signal Y_1, Y_1_d1 :  std_logic_vector(24 downto 0);
   -- timing of Y_1: (c2, 1.180000ns)
signal S_1 :  std_logic_vector(24 downto 0);
   -- timing of S_1: (c3, 0.620000ns)
signal R_1 :  std_logic_vector(23 downto 0);
   -- timing of R_1: (c3, 0.620000ns)
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            Cin_1_d1 <=  Cin_1;
            Cin_1_d2 <=  Cin_1_d1;
            Cin_1_d3 <=  Cin_1_d2;
            X_1_d1 <=  X_1;
            Y_1_d1 <=  Y_1;
         end if;
      end process;
   Cin_1 <= Cin;
   X_1 <= '0' & X(23 downto 0);
   Y_1 <= '0' & Y(23 downto 0);
   S_1 <= X_1_d1 + Y_1_d1 + Cin_1_d3;
   R_1 <= S_1(23 downto 0);
   R <= R_1 ;
end architecture;

--------------------------------------------------------------------------------
--                         IntAdder_24_Freq500_uid25
-- VHDL generated for DummyFPGA @ 500MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin (2008-2016)
--------------------------------------------------------------------------------
-- Pipeline depth: 6 cycles
-- Clock period (ns): 2
-- Target frequency (MHz): 500
-- Input signals: X Y Cin
-- Output signals: R
--  approx. input signal timings: X: (c3, 0.620000ns)Y: (c5, 0.675385ns)Cin: (c0, 0.000000ns)
--  approx. output signal timings: R: (c6, 0.105385ns)

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntAdder_24_Freq500_uid25 is
    port (clk : in std_logic;
          X : in  std_logic_vector(23 downto 0);
          Y : in  std_logic_vector(23 downto 0);
          Cin : in  std_logic;
          R : out  std_logic_vector(23 downto 0)   );
end entity;

architecture arch of IntAdder_24_Freq500_uid25 is
signal Rtmp :  std_logic_vector(23 downto 0);
   -- timing of Rtmp: (c6, 0.105385ns)
signal X_d1, X_d2, X_d3 :  std_logic_vector(23 downto 0);
   -- timing of X: (c3, 0.620000ns)
signal Y_d1 :  std_logic_vector(23 downto 0);
   -- timing of Y: (c5, 0.675385ns)
signal Cin_d1, Cin_d2, Cin_d3, Cin_d4, Cin_d5, Cin_d6 :  std_logic;
   -- timing of Cin: (c0, 0.000000ns)
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            X_d1 <=  X;
            X_d2 <=  X_d1;
            X_d3 <=  X_d2;
            Y_d1 <=  Y;
            Cin_d1 <=  Cin;
            Cin_d2 <=  Cin_d1;
            Cin_d3 <=  Cin_d2;
            Cin_d4 <=  Cin_d3;
            Cin_d5 <=  Cin_d4;
            Cin_d6 <=  Cin_d5;
         end if;
      end process;
   Rtmp <= X_d3 + Y_d1 + Cin_d6;
   R <= Rtmp;
end architecture;

--------------------------------------------------------------------------------
--                         IntAdder_35_Freq500_uid34
-- VHDL generated for DummyFPGA @ 500MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin (2008-2016)
--------------------------------------------------------------------------------
-- Pipeline depth: 2 cycles
-- Clock period (ns): 2
-- Target frequency (MHz): 500
-- Input signals: X Y Cin
-- Output signals: R
--  approx. input signal timings: X: (c0, 0.550000ns)Y: (c1, 1.200000ns)Cin: (c0, 0.000000ns)
--  approx. output signal timings: R: (c2, 0.750000ns)

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntAdder_35_Freq500_uid34 is
    port (clk : in std_logic;
          X : in  std_logic_vector(34 downto 0);
          Y : in  std_logic_vector(34 downto 0);
          Cin : in  std_logic;
          R : out  std_logic_vector(34 downto 0)   );
end entity;

architecture arch of IntAdder_35_Freq500_uid34 is
signal Cin_1, Cin_1_d1, Cin_1_d2 :  std_logic;
   -- timing of Cin_1: (c0, 0.000000ns)
signal X_1, X_1_d1, X_1_d2 :  std_logic_vector(35 downto 0);
   -- timing of X_1: (c0, 0.550000ns)
signal Y_1, Y_1_d1 :  std_logic_vector(35 downto 0);
   -- timing of Y_1: (c1, 1.200000ns)
signal S_1 :  std_logic_vector(35 downto 0);
   -- timing of S_1: (c2, 0.750000ns)
signal R_1 :  std_logic_vector(34 downto 0);
   -- timing of R_1: (c2, 0.750000ns)
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            Cin_1_d1 <=  Cin_1;
            Cin_1_d2 <=  Cin_1_d1;
            X_1_d1 <=  X_1;
            X_1_d2 <=  X_1_d1;
            Y_1_d1 <=  Y_1;
         end if;
      end process;
   Cin_1 <= Cin;
   X_1 <= '0' & X(34 downto 0);
   Y_1 <= '0' & Y(34 downto 0);
   S_1 <= X_1_d2 + Y_1_d1 + Cin_1_d2;
   R_1 <= S_1(34 downto 0);
   R <= R_1 ;
end architecture;

--------------------------------------------------------------------------------
--                         IntAdder_35_Freq500_uid37
-- VHDL generated for DummyFPGA @ 500MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin (2008-2016)
--------------------------------------------------------------------------------
-- Pipeline depth: 6 cycles
-- Clock period (ns): 2
-- Target frequency (MHz): 500
-- Input signals: X Y Cin
-- Output signals: R
--  approx. input signal timings: X: (c2, 0.750000ns)Y: (c6, 0.105385ns)Cin: (c0, 0.000000ns)
--  approx. output signal timings: R: (c6, 1.445385ns)

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntAdder_35_Freq500_uid37 is
    port (clk : in std_logic;
          X : in  std_logic_vector(34 downto 0);
          Y : in  std_logic_vector(34 downto 0);
          Cin : in  std_logic;
          R : out  std_logic_vector(34 downto 0)   );
end entity;

architecture arch of IntAdder_35_Freq500_uid37 is
signal Rtmp :  std_logic_vector(34 downto 0);
   -- timing of Rtmp: (c6, 1.445385ns)
signal X_d1, X_d2, X_d3, X_d4 :  std_logic_vector(34 downto 0);
   -- timing of X: (c2, 0.750000ns)
signal Cin_d1, Cin_d2, Cin_d3, Cin_d4, Cin_d5, Cin_d6 :  std_logic;
   -- timing of Cin: (c0, 0.000000ns)
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            X_d1 <=  X;
            X_d2 <=  X_d1;
            X_d3 <=  X_d2;
            X_d4 <=  X_d3;
            Cin_d1 <=  Cin;
            Cin_d2 <=  Cin_d1;
            Cin_d3 <=  Cin_d2;
            Cin_d4 <=  Cin_d3;
            Cin_d5 <=  Cin_d4;
            Cin_d6 <=  Cin_d5;
         end if;
      end process;
   Rtmp <= X_d4 + Y + Cin_d6;
   R <= Rtmp;
end architecture;

--------------------------------------------------------------------------------
--                         IntAdder_32_Freq500_uid49
-- VHDL generated for DummyFPGA @ 500MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin (2008-2016)
--------------------------------------------------------------------------------
-- Pipeline depth: 1 cycles
-- Clock period (ns): 2
-- Target frequency (MHz): 500
-- Input signals: X Y Cin
-- Output signals: R
--  approx. input signal timings: X: (c1, 0.370000ns)Y: (c1, 0.370000ns)Cin: (c0, 0.000000ns)
--  approx. output signal timings: R: (c1, 1.680000ns)

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntAdder_32_Freq500_uid49 is
    port (clk : in std_logic;
          X : in  std_logic_vector(31 downto 0);
          Y : in  std_logic_vector(31 downto 0);
          Cin : in  std_logic;
          R : out  std_logic_vector(31 downto 0)   );
end entity;

architecture arch of IntAdder_32_Freq500_uid49 is
signal Rtmp :  std_logic_vector(31 downto 0);
   -- timing of Rtmp: (c1, 1.680000ns)
signal Cin_d1 :  std_logic;
   -- timing of Cin: (c0, 0.000000ns)
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            Cin_d1 <=  Cin;
         end if;
      end process;
   Rtmp <= X + Y + Cin_d1;
   R <= Rtmp;
end architecture;

--------------------------------------------------------------------------------
--                          FixRealKCM_Freq500_uid39
-- VHDL generated for DummyFPGA @ 500MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin (2007-2016)
--------------------------------------------------------------------------------
-- Pipeline depth: 1 cycles
-- Clock period (ns): 2
-- Target frequency (MHz): 500
-- Input signals: X
-- Output signals: R
--  approx. input signal timings: X: (c0, 1.620000ns)
--  approx. output signal timings: R: (c1, 1.680000ns)

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity FixRealKCM_Freq500_uid39 is
    port (clk : in std_logic;
          X : in  std_logic_vector(7 downto 0);
          R : out  std_logic_vector(31 downto 0)   );
end entity;

architecture arch of FixRealKCM_Freq500_uid39 is
   component FixRealKCM_Freq500_uid39_T0_Freq500_uid42 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(31 downto 0)   );
   end component;

   component FixRealKCM_Freq500_uid39_T1_Freq500_uid45 is
      port ( X : in  std_logic_vector(2 downto 0);
             Y : out  std_logic_vector(26 downto 0)   );
   end component;

   component IntAdder_32_Freq500_uid49 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(31 downto 0);
             Y : in  std_logic_vector(31 downto 0);
             Cin : in  std_logic;
             R : out  std_logic_vector(31 downto 0)   );
   end component;

signal FixRealKCM_Freq500_uid39_A0 :  std_logic_vector(4 downto 0);
   -- timing of FixRealKCM_Freq500_uid39_A0: (c0, 1.620000ns)
signal FixRealKCM_Freq500_uid39_T0 :  std_logic_vector(31 downto 0);
   -- timing of FixRealKCM_Freq500_uid39_T0: (c1, 0.370000ns)
signal FixRealKCM_Freq500_uid39_T0_copy43, FixRealKCM_Freq500_uid39_T0_copy43_d1 :  std_logic_vector(31 downto 0);
   -- timing of FixRealKCM_Freq500_uid39_T0_copy43: (c0, 1.620000ns)
signal bh40_w0_0 :  std_logic;
   -- timing of bh40_w0_0: (c1, 0.370000ns)
signal bh40_w1_0 :  std_logic;
   -- timing of bh40_w1_0: (c1, 0.370000ns)
signal bh40_w2_0 :  std_logic;
   -- timing of bh40_w2_0: (c1, 0.370000ns)
signal bh40_w3_0 :  std_logic;
   -- timing of bh40_w3_0: (c1, 0.370000ns)
signal bh40_w4_0 :  std_logic;
   -- timing of bh40_w4_0: (c1, 0.370000ns)
signal bh40_w5_0 :  std_logic;
   -- timing of bh40_w5_0: (c1, 0.370000ns)
signal bh40_w6_0 :  std_logic;
   -- timing of bh40_w6_0: (c1, 0.370000ns)
signal bh40_w7_0 :  std_logic;
   -- timing of bh40_w7_0: (c1, 0.370000ns)
signal bh40_w8_0 :  std_logic;
   -- timing of bh40_w8_0: (c1, 0.370000ns)
signal bh40_w9_0 :  std_logic;
   -- timing of bh40_w9_0: (c1, 0.370000ns)
signal bh40_w10_0 :  std_logic;
   -- timing of bh40_w10_0: (c1, 0.370000ns)
signal bh40_w11_0 :  std_logic;
   -- timing of bh40_w11_0: (c1, 0.370000ns)
signal bh40_w12_0 :  std_logic;
   -- timing of bh40_w12_0: (c1, 0.370000ns)
signal bh40_w13_0 :  std_logic;
   -- timing of bh40_w13_0: (c1, 0.370000ns)
signal bh40_w14_0 :  std_logic;
   -- timing of bh40_w14_0: (c1, 0.370000ns)
signal bh40_w15_0 :  std_logic;
   -- timing of bh40_w15_0: (c1, 0.370000ns)
signal bh40_w16_0 :  std_logic;
   -- timing of bh40_w16_0: (c1, 0.370000ns)
signal bh40_w17_0 :  std_logic;
   -- timing of bh40_w17_0: (c1, 0.370000ns)
signal bh40_w18_0 :  std_logic;
   -- timing of bh40_w18_0: (c1, 0.370000ns)
signal bh40_w19_0 :  std_logic;
   -- timing of bh40_w19_0: (c1, 0.370000ns)
signal bh40_w20_0 :  std_logic;
   -- timing of bh40_w20_0: (c1, 0.370000ns)
signal bh40_w21_0 :  std_logic;
   -- timing of bh40_w21_0: (c1, 0.370000ns)
signal bh40_w22_0 :  std_logic;
   -- timing of bh40_w22_0: (c1, 0.370000ns)
signal bh40_w23_0 :  std_logic;
   -- timing of bh40_w23_0: (c1, 0.370000ns)
signal bh40_w24_0 :  std_logic;
   -- timing of bh40_w24_0: (c1, 0.370000ns)
signal bh40_w25_0 :  std_logic;
   -- timing of bh40_w25_0: (c1, 0.370000ns)
signal bh40_w26_0 :  std_logic;
   -- timing of bh40_w26_0: (c1, 0.370000ns)
signal bh40_w27_0 :  std_logic;
   -- timing of bh40_w27_0: (c1, 0.370000ns)
signal bh40_w28_0 :  std_logic;
   -- timing of bh40_w28_0: (c1, 0.370000ns)
signal bh40_w29_0 :  std_logic;
   -- timing of bh40_w29_0: (c1, 0.370000ns)
signal bh40_w30_0 :  std_logic;
   -- timing of bh40_w30_0: (c1, 0.370000ns)
signal bh40_w31_0 :  std_logic;
   -- timing of bh40_w31_0: (c1, 0.370000ns)
signal FixRealKCM_Freq500_uid39_A1 :  std_logic_vector(2 downto 0);
   -- timing of FixRealKCM_Freq500_uid39_A1: (c0, 1.620000ns)
signal FixRealKCM_Freq500_uid39_T1 :  std_logic_vector(26 downto 0);
   -- timing of FixRealKCM_Freq500_uid39_T1: (c1, 0.370000ns)
signal FixRealKCM_Freq500_uid39_T1_copy46, FixRealKCM_Freq500_uid39_T1_copy46_d1 :  std_logic_vector(26 downto 0);
   -- timing of FixRealKCM_Freq500_uid39_T1_copy46: (c0, 1.620000ns)
signal bh40_w0_1 :  std_logic;
   -- timing of bh40_w0_1: (c1, 0.370000ns)
signal bh40_w1_1 :  std_logic;
   -- timing of bh40_w1_1: (c1, 0.370000ns)
signal bh40_w2_1 :  std_logic;
   -- timing of bh40_w2_1: (c1, 0.370000ns)
signal bh40_w3_1 :  std_logic;
   -- timing of bh40_w3_1: (c1, 0.370000ns)
signal bh40_w4_1 :  std_logic;
   -- timing of bh40_w4_1: (c1, 0.370000ns)
signal bh40_w5_1 :  std_logic;
   -- timing of bh40_w5_1: (c1, 0.370000ns)
signal bh40_w6_1 :  std_logic;
   -- timing of bh40_w6_1: (c1, 0.370000ns)
signal bh40_w7_1 :  std_logic;
   -- timing of bh40_w7_1: (c1, 0.370000ns)
signal bh40_w8_1 :  std_logic;
   -- timing of bh40_w8_1: (c1, 0.370000ns)
signal bh40_w9_1 :  std_logic;
   -- timing of bh40_w9_1: (c1, 0.370000ns)
signal bh40_w10_1 :  std_logic;
   -- timing of bh40_w10_1: (c1, 0.370000ns)
signal bh40_w11_1 :  std_logic;
   -- timing of bh40_w11_1: (c1, 0.370000ns)
signal bh40_w12_1 :  std_logic;
   -- timing of bh40_w12_1: (c1, 0.370000ns)
signal bh40_w13_1 :  std_logic;
   -- timing of bh40_w13_1: (c1, 0.370000ns)
signal bh40_w14_1 :  std_logic;
   -- timing of bh40_w14_1: (c1, 0.370000ns)
signal bh40_w15_1 :  std_logic;
   -- timing of bh40_w15_1: (c1, 0.370000ns)
signal bh40_w16_1 :  std_logic;
   -- timing of bh40_w16_1: (c1, 0.370000ns)
signal bh40_w17_1 :  std_logic;
   -- timing of bh40_w17_1: (c1, 0.370000ns)
signal bh40_w18_1 :  std_logic;
   -- timing of bh40_w18_1: (c1, 0.370000ns)
signal bh40_w19_1 :  std_logic;
   -- timing of bh40_w19_1: (c1, 0.370000ns)
signal bh40_w20_1 :  std_logic;
   -- timing of bh40_w20_1: (c1, 0.370000ns)
signal bh40_w21_1 :  std_logic;
   -- timing of bh40_w21_1: (c1, 0.370000ns)
signal bh40_w22_1 :  std_logic;
   -- timing of bh40_w22_1: (c1, 0.370000ns)
signal bh40_w23_1 :  std_logic;
   -- timing of bh40_w23_1: (c1, 0.370000ns)
signal bh40_w24_1 :  std_logic;
   -- timing of bh40_w24_1: (c1, 0.370000ns)
signal bh40_w25_1 :  std_logic;
   -- timing of bh40_w25_1: (c1, 0.370000ns)
signal bh40_w26_1 :  std_logic;
   -- timing of bh40_w26_1: (c1, 0.370000ns)
signal bitheapFinalAdd_bh40_In0 :  std_logic_vector(31 downto 0);
   -- timing of bitheapFinalAdd_bh40_In0: (c1, 0.370000ns)
signal bitheapFinalAdd_bh40_In1 :  std_logic_vector(31 downto 0);
   -- timing of bitheapFinalAdd_bh40_In1: (c1, 0.370000ns)
signal bitheapFinalAdd_bh40_Cin :  std_logic;
   -- timing of bitheapFinalAdd_bh40_Cin: (c0, 0.000000ns)
signal bitheapFinalAdd_bh40_Out :  std_logic_vector(31 downto 0);
   -- timing of bitheapFinalAdd_bh40_Out: (c1, 1.680000ns)
signal bitheapResult_bh40 :  std_logic_vector(31 downto 0);
   -- timing of bitheapResult_bh40: (c1, 1.680000ns)
signal OutRes :  std_logic_vector(31 downto 0);
   -- timing of OutRes: (c1, 1.680000ns)
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            FixRealKCM_Freq500_uid39_T0_copy43_d1 <=  FixRealKCM_Freq500_uid39_T0_copy43;
            FixRealKCM_Freq500_uid39_T1_copy46_d1 <=  FixRealKCM_Freq500_uid39_T1_copy46;
         end if;
      end process;
-- This operator multiplies by log(2)
   FixRealKCM_Freq500_uid39_A0 <= X(7 downto 3);-- input address  m=7  l=3
   FixRealKCM_Freq500_uid39_Table0: FixRealKCM_Freq500_uid39_T0_Freq500_uid42
      port map ( X => FixRealKCM_Freq500_uid39_A0,
                 Y => FixRealKCM_Freq500_uid39_T0_copy43);
   FixRealKCM_Freq500_uid39_T0 <= FixRealKCM_Freq500_uid39_T0_copy43_d1; -- output copy to hold a pipeline register if needed
   bh40_w0_0 <= FixRealKCM_Freq500_uid39_T0(0);
   bh40_w1_0 <= FixRealKCM_Freq500_uid39_T0(1);
   bh40_w2_0 <= FixRealKCM_Freq500_uid39_T0(2);
   bh40_w3_0 <= FixRealKCM_Freq500_uid39_T0(3);
   bh40_w4_0 <= FixRealKCM_Freq500_uid39_T0(4);
   bh40_w5_0 <= FixRealKCM_Freq500_uid39_T0(5);
   bh40_w6_0 <= FixRealKCM_Freq500_uid39_T0(6);
   bh40_w7_0 <= FixRealKCM_Freq500_uid39_T0(7);
   bh40_w8_0 <= FixRealKCM_Freq500_uid39_T0(8);
   bh40_w9_0 <= FixRealKCM_Freq500_uid39_T0(9);
   bh40_w10_0 <= FixRealKCM_Freq500_uid39_T0(10);
   bh40_w11_0 <= FixRealKCM_Freq500_uid39_T0(11);
   bh40_w12_0 <= FixRealKCM_Freq500_uid39_T0(12);
   bh40_w13_0 <= FixRealKCM_Freq500_uid39_T0(13);
   bh40_w14_0 <= FixRealKCM_Freq500_uid39_T0(14);
   bh40_w15_0 <= FixRealKCM_Freq500_uid39_T0(15);
   bh40_w16_0 <= FixRealKCM_Freq500_uid39_T0(16);
   bh40_w17_0 <= FixRealKCM_Freq500_uid39_T0(17);
   bh40_w18_0 <= FixRealKCM_Freq500_uid39_T0(18);
   bh40_w19_0 <= FixRealKCM_Freq500_uid39_T0(19);
   bh40_w20_0 <= FixRealKCM_Freq500_uid39_T0(20);
   bh40_w21_0 <= FixRealKCM_Freq500_uid39_T0(21);
   bh40_w22_0 <= FixRealKCM_Freq500_uid39_T0(22);
   bh40_w23_0 <= FixRealKCM_Freq500_uid39_T0(23);
   bh40_w24_0 <= FixRealKCM_Freq500_uid39_T0(24);
   bh40_w25_0 <= FixRealKCM_Freq500_uid39_T0(25);
   bh40_w26_0 <= FixRealKCM_Freq500_uid39_T0(26);
   bh40_w27_0 <= FixRealKCM_Freq500_uid39_T0(27);
   bh40_w28_0 <= FixRealKCM_Freq500_uid39_T0(28);
   bh40_w29_0 <= FixRealKCM_Freq500_uid39_T0(29);
   bh40_w30_0 <= FixRealKCM_Freq500_uid39_T0(30);
   bh40_w31_0 <= FixRealKCM_Freq500_uid39_T0(31);
   FixRealKCM_Freq500_uid39_A1 <= X(2 downto 0);-- input address  m=2  l=0
   FixRealKCM_Freq500_uid39_Table1: FixRealKCM_Freq500_uid39_T1_Freq500_uid45
      port map ( X => FixRealKCM_Freq500_uid39_A1,
                 Y => FixRealKCM_Freq500_uid39_T1_copy46);
   FixRealKCM_Freq500_uid39_T1 <= FixRealKCM_Freq500_uid39_T1_copy46_d1; -- output copy to hold a pipeline register if needed
   bh40_w0_1 <= FixRealKCM_Freq500_uid39_T1(0);
   bh40_w1_1 <= FixRealKCM_Freq500_uid39_T1(1);
   bh40_w2_1 <= FixRealKCM_Freq500_uid39_T1(2);
   bh40_w3_1 <= FixRealKCM_Freq500_uid39_T1(3);
   bh40_w4_1 <= FixRealKCM_Freq500_uid39_T1(4);
   bh40_w5_1 <= FixRealKCM_Freq500_uid39_T1(5);
   bh40_w6_1 <= FixRealKCM_Freq500_uid39_T1(6);
   bh40_w7_1 <= FixRealKCM_Freq500_uid39_T1(7);
   bh40_w8_1 <= FixRealKCM_Freq500_uid39_T1(8);
   bh40_w9_1 <= FixRealKCM_Freq500_uid39_T1(9);
   bh40_w10_1 <= FixRealKCM_Freq500_uid39_T1(10);
   bh40_w11_1 <= FixRealKCM_Freq500_uid39_T1(11);
   bh40_w12_1 <= FixRealKCM_Freq500_uid39_T1(12);
   bh40_w13_1 <= FixRealKCM_Freq500_uid39_T1(13);
   bh40_w14_1 <= FixRealKCM_Freq500_uid39_T1(14);
   bh40_w15_1 <= FixRealKCM_Freq500_uid39_T1(15);
   bh40_w16_1 <= FixRealKCM_Freq500_uid39_T1(16);
   bh40_w17_1 <= FixRealKCM_Freq500_uid39_T1(17);
   bh40_w18_1 <= FixRealKCM_Freq500_uid39_T1(18);
   bh40_w19_1 <= FixRealKCM_Freq500_uid39_T1(19);
   bh40_w20_1 <= FixRealKCM_Freq500_uid39_T1(20);
   bh40_w21_1 <= FixRealKCM_Freq500_uid39_T1(21);
   bh40_w22_1 <= FixRealKCM_Freq500_uid39_T1(22);
   bh40_w23_1 <= FixRealKCM_Freq500_uid39_T1(23);
   bh40_w24_1 <= FixRealKCM_Freq500_uid39_T1(24);
   bh40_w25_1 <= FixRealKCM_Freq500_uid39_T1(25);
   bh40_w26_1 <= FixRealKCM_Freq500_uid39_T1(26);

   -- Adding the constant bits 
      -- All the constant bits are zero, nothing to add


   bitheapFinalAdd_bh40_In0 <= "" & bh40_w31_0 & bh40_w30_0 & bh40_w29_0 & bh40_w28_0 & bh40_w27_0 & bh40_w26_1 & bh40_w25_1 & bh40_w24_1 & bh40_w23_1 & bh40_w22_1 & bh40_w21_1 & bh40_w20_1 & bh40_w19_1 & bh40_w18_1 & bh40_w17_1 & bh40_w16_1 & bh40_w15_1 & bh40_w14_1 & bh40_w13_1 & bh40_w12_1 & bh40_w11_1 & bh40_w10_1 & bh40_w9_1 & bh40_w8_1 & bh40_w7_1 & bh40_w6_1 & bh40_w5_1 & bh40_w4_1 & bh40_w3_1 & bh40_w2_1 & bh40_w1_1 & bh40_w0_1;
   bitheapFinalAdd_bh40_In1 <= "0" & "0" & "0" & "0" & "0" & bh40_w26_0 & bh40_w25_0 & bh40_w24_0 & bh40_w23_0 & bh40_w22_0 & bh40_w21_0 & bh40_w20_0 & bh40_w19_0 & bh40_w18_0 & bh40_w17_0 & bh40_w16_0 & bh40_w15_0 & bh40_w14_0 & bh40_w13_0 & bh40_w12_0 & bh40_w11_0 & bh40_w10_0 & bh40_w9_0 & bh40_w8_0 & bh40_w7_0 & bh40_w6_0 & bh40_w5_0 & bh40_w4_0 & bh40_w3_0 & bh40_w2_0 & bh40_w1_0 & bh40_w0_0;
   bitheapFinalAdd_bh40_Cin <= '0';

   bitheapFinalAdd_bh40: IntAdder_32_Freq500_uid49
      port map ( clk  => clk,
                 Cin => bitheapFinalAdd_bh40_Cin,
                 X => bitheapFinalAdd_bh40_In0,
                 Y => bitheapFinalAdd_bh40_In1,
                 R => bitheapFinalAdd_bh40_Out);
   bitheapResult_bh40 <= bitheapFinalAdd_bh40_Out(31 downto 0);
   OutRes <= bitheapResult_bh40(31 downto 0);
   R <= OutRes(31 downto 0);
end architecture;

--------------------------------------------------------------------------------
--                         IntAdder_43_Freq500_uid51
-- VHDL generated for DummyFPGA @ 500MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin (2008-2016)
--------------------------------------------------------------------------------
-- Pipeline depth: 8 cycles
-- Clock period (ns): 2
-- Target frequency (MHz): 500
-- Input signals: X Y Cin
-- Output signals: R
--  approx. input signal timings: X: (c1, 1.680000ns)Y: (c6, 1.445385ns)Cin: (c0, 0.550000ns)
--  approx. output signal timings: R: (c8, 0.275385ns)

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntAdder_43_Freq500_uid51 is
    port (clk : in std_logic;
          X : in  std_logic_vector(42 downto 0);
          Y : in  std_logic_vector(42 downto 0);
          Cin : in  std_logic;
          R : out  std_logic_vector(42 downto 0)   );
end entity;

architecture arch of IntAdder_43_Freq500_uid51 is
signal Cin_0, Cin_0_d1, Cin_0_d2, Cin_0_d3, Cin_0_d4, Cin_0_d5, Cin_0_d6, Cin_0_d7 :  std_logic;
   -- timing of Cin_0: (c0, 0.550000ns)
signal X_0, X_0_d1, X_0_d2, X_0_d3, X_0_d4, X_0_d5, X_0_d6 :  std_logic_vector(25 downto 0);
   -- timing of X_0: (c1, 1.680000ns)
signal Y_0, Y_0_d1 :  std_logic_vector(25 downto 0);
   -- timing of Y_0: (c6, 1.445385ns)
signal S_0 :  std_logic_vector(25 downto 0);
   -- timing of S_0: (c7, 0.895385ns)
signal R_0, R_0_d1 :  std_logic_vector(24 downto 0);
   -- timing of R_0: (c7, 0.895385ns)
signal Cin_1, Cin_1_d1 :  std_logic;
   -- timing of Cin_1: (c7, 0.895385ns)
signal X_1, X_1_d1, X_1_d2, X_1_d3, X_1_d4, X_1_d5, X_1_d6, X_1_d7 :  std_logic_vector(18 downto 0);
   -- timing of X_1: (c1, 1.680000ns)
signal Y_1, Y_1_d1, Y_1_d2 :  std_logic_vector(18 downto 0);
   -- timing of Y_1: (c6, 1.445385ns)
signal S_1 :  std_logic_vector(18 downto 0);
   -- timing of S_1: (c8, 0.275385ns)
signal R_1 :  std_logic_vector(17 downto 0);
   -- timing of R_1: (c8, 0.275385ns)
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            Cin_0_d1 <=  Cin_0;
            Cin_0_d2 <=  Cin_0_d1;
            Cin_0_d3 <=  Cin_0_d2;
            Cin_0_d4 <=  Cin_0_d3;
            Cin_0_d5 <=  Cin_0_d4;
            Cin_0_d6 <=  Cin_0_d5;
            Cin_0_d7 <=  Cin_0_d6;
            X_0_d1 <=  X_0;
            X_0_d2 <=  X_0_d1;
            X_0_d3 <=  X_0_d2;
            X_0_d4 <=  X_0_d3;
            X_0_d5 <=  X_0_d4;
            X_0_d6 <=  X_0_d5;
            Y_0_d1 <=  Y_0;
            R_0_d1 <=  R_0;
            Cin_1_d1 <=  Cin_1;
            X_1_d1 <=  X_1;
            X_1_d2 <=  X_1_d1;
            X_1_d3 <=  X_1_d2;
            X_1_d4 <=  X_1_d3;
            X_1_d5 <=  X_1_d4;
            X_1_d6 <=  X_1_d5;
            X_1_d7 <=  X_1_d6;
            Y_1_d1 <=  Y_1;
            Y_1_d2 <=  Y_1_d1;
         end if;
      end process;
   Cin_0 <= Cin;
   X_0 <= '0' & X(24 downto 0);
   Y_0 <= '0' & Y(24 downto 0);
   S_0 <= X_0_d6 + Y_0_d1 + Cin_0_d7;
   R_0 <= S_0(24 downto 0);
   Cin_1 <= S_0(25);
   X_1 <= '0' & X(42 downto 25);
   Y_1 <= '0' & Y(42 downto 25);
   S_1 <= X_1_d7 + Y_1_d2 + Cin_1_d1;
   R_1 <= S_1(17 downto 0);
   R <= R_1 & R_0_d1 ;
end architecture;

--------------------------------------------------------------------------------
--                    Normalizer_Z_43_35_18_Freq500_uid53
-- VHDL generated for DummyFPGA @ 500MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, (2007-2020)
--------------------------------------------------------------------------------
-- Pipeline depth: 3 cycles
-- Clock period (ns): 2
-- Target frequency (MHz): 500
-- Input signals: X
-- Output signals: Count R
--  approx. input signal timings: X: (c8, 0.275385ns)
--  approx. output signal timings: Count: (c10, 1.715385ns)R: (c11, 0.465385ns)

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity Normalizer_Z_43_35_18_Freq500_uid53 is
    port (clk : in std_logic;
          X : in  std_logic_vector(42 downto 0);
          Count : out  std_logic_vector(4 downto 0);
          R : out  std_logic_vector(34 downto 0)   );
end entity;

architecture arch of Normalizer_Z_43_35_18_Freq500_uid53 is
signal level5 :  std_logic_vector(42 downto 0);
   -- timing of level5: (c8, 0.275385ns)
signal count4, count4_d1, count4_d2 :  std_logic;
   -- timing of count4: (c8, 0.865385ns)
signal level4, level4_d1 :  std_logic_vector(42 downto 0);
   -- timing of level4: (c8, 1.415385ns)
signal count3, count3_d1 :  std_logic;
   -- timing of count3: (c9, 0.185385ns)
signal level3, level3_d1 :  std_logic_vector(41 downto 0);
   -- timing of level3: (c9, 0.735385ns)
signal count2, count2_d1 :  std_logic;
   -- timing of count2: (c9, 1.295385ns)
signal level2 :  std_logic_vector(37 downto 0);
   -- timing of level2: (c10, 0.045385ns)
signal count1 :  std_logic;
   -- timing of count1: (c10, 0.605385ns)
signal level1, level1_d1 :  std_logic_vector(35 downto 0);
   -- timing of level1: (c10, 1.155385ns)
signal count0, count0_d1 :  std_logic;
   -- timing of count0: (c10, 1.715385ns)
signal level0 :  std_logic_vector(34 downto 0);
   -- timing of level0: (c11, 0.465385ns)
signal sCount :  std_logic_vector(4 downto 0);
   -- timing of sCount: (c10, 1.715385ns)
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            count4_d1 <=  count4;
            count4_d2 <=  count4_d1;
            level4_d1 <=  level4;
            count3_d1 <=  count3;
            level3_d1 <=  level3;
            count2_d1 <=  count2;
            level1_d1 <=  level1;
            count0_d1 <=  count0;
         end if;
      end process;
   level5 <= X ;
   count4<= '1' when level5(42 downto 27) = (42 downto 27=>'0') else '0';
   level4<= level5(42 downto 0) when count4='0' else level5(26 downto 0) & (15 downto 0 => '0');

   count3<= '1' when level4_d1(42 downto 35) = (42 downto 35=>'0') else '0';
   level3<= level4_d1(42 downto 1) when count3='0' else level4_d1(34 downto 0) & (6 downto 0 => '0');

   count2<= '1' when level3(41 downto 38) = (41 downto 38=>'0') else '0';
   level2<= level3_d1(41 downto 4) when count2_d1='0' else level3_d1(37 downto 0);

   count1<= '1' when level2(37 downto 36) = (37 downto 36=>'0') else '0';
   level1<= level2(37 downto 2) when count1='0' else level2(35 downto 0);

   count0<= '1' when level1(35 downto 35) = (35 downto 35=>'0') else '0';
   level0<= level1_d1(35 downto 1) when count0_d1='0' else level1_d1(34 downto 0);

   R <= level0;
   sCount <= count4_d2 & count3_d1 & count2_d1 & count1 & count0;
   Count <= sCount;
end architecture;

--------------------------------------------------------------------------------
--                   RightShifter15_by_max_14_Freq500_uid55
-- VHDL generated for DummyFPGA @ 500MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca (2008-2011), Florent de Dinechin (2008-2019)
--------------------------------------------------------------------------------
-- Pipeline depth: 3 cycles
-- Clock period (ns): 2
-- Target frequency (MHz): 500
-- Input signals: X S
-- Output signals: R
--  approx. input signal timings: X: (c5, 0.125385ns)S: (c3, 1.460000ns)
--  approx. output signal timings: R: (c6, 0.163846ns)

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity RightShifter15_by_max_14_Freq500_uid55 is
    port (clk : in std_logic;
          X : in  std_logic_vector(14 downto 0);
          S : in  std_logic_vector(3 downto 0);
          R : out  std_logic_vector(28 downto 0)   );
end entity;

architecture arch of RightShifter15_by_max_14_Freq500_uid55 is
signal ps, ps_d1, ps_d2, ps_d3 :  std_logic_vector(3 downto 0);
   -- timing of ps: (c3, 1.460000ns)
signal level0 :  std_logic_vector(14 downto 0);
   -- timing of level0: (c5, 0.125385ns)
signal level1 :  std_logic_vector(15 downto 0);
   -- timing of level1: (c5, 0.125385ns)
signal level2 :  std_logic_vector(17 downto 0);
   -- timing of level2: (c5, 0.952308ns)
signal level3, level3_d1 :  std_logic_vector(21 downto 0);
   -- timing of level3: (c5, 0.952308ns)
signal level4 :  std_logic_vector(29 downto 0);
   -- timing of level4: (c6, 0.163846ns)
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            ps_d1 <=  ps;
            ps_d2 <=  ps_d1;
            ps_d3 <=  ps_d2;
            level3_d1 <=  level3;
         end if;
      end process;
   ps<= S;
   level0<= X;
   level1 <=  (0 downto 0 => '0') & level0 when ps_d2(0) = '1' else    level0 & (0 downto 0 => '0');
   level2 <=  (1 downto 0 => '0') & level1 when ps_d2(1) = '1' else    level1 & (1 downto 0 => '0');
   level3 <=  (3 downto 0 => '0') & level2 when ps_d2(2) = '1' else    level2 & (3 downto 0 => '0');
   level4 <=  (7 downto 0 => '0') & level3_d1 when ps_d3(3) = '1' else    level3_d1 & (7 downto 0 => '0');
   R <= level4(29 downto 1);
end architecture;

--------------------------------------------------------------------------------
--                         IntAdder_26_Freq500_uid57
-- VHDL generated for DummyFPGA @ 500MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin (2008-2016)
--------------------------------------------------------------------------------
-- Pipeline depth: 6 cycles
-- Clock period (ns): 2
-- Target frequency (MHz): 500
-- Input signals: X Y Cin
-- Output signals: R
--  approx. input signal timings: X: (c4, 1.375385ns)Y: (c6, 0.163846ns)Cin: (c0, 0.550000ns)
--  approx. output signal timings: R: (c6, 1.413846ns)

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntAdder_26_Freq500_uid57 is
    port (clk : in std_logic;
          X : in  std_logic_vector(25 downto 0);
          Y : in  std_logic_vector(25 downto 0);
          Cin : in  std_logic;
          R : out  std_logic_vector(25 downto 0)   );
end entity;

architecture arch of IntAdder_26_Freq500_uid57 is
signal Rtmp :  std_logic_vector(25 downto 0);
   -- timing of Rtmp: (c6, 1.413846ns)
signal X_d1, X_d2 :  std_logic_vector(25 downto 0);
   -- timing of X: (c4, 1.375385ns)
signal Cin_d1, Cin_d2, Cin_d3, Cin_d4, Cin_d5, Cin_d6 :  std_logic;
   -- timing of Cin: (c0, 0.550000ns)
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            X_d1 <=  X;
            X_d2 <=  X_d1;
            Cin_d1 <=  Cin;
            Cin_d2 <=  Cin_d1;
            Cin_d3 <=  Cin_d2;
            Cin_d4 <=  Cin_d3;
            Cin_d5 <=  Cin_d4;
            Cin_d6 <=  Cin_d5;
         end if;
      end process;
   Rtmp <= X_d2 + Y + Cin_d6;
   R <= Rtmp;
end architecture;

--------------------------------------------------------------------------------
--                         IntAdder_28_Freq500_uid60
-- VHDL generated for DummyFPGA @ 500MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin (2008-2016)
--------------------------------------------------------------------------------
-- Pipeline depth: 11 cycles
-- Clock period (ns): 2
-- Target frequency (MHz): 500
-- Input signals: X Y Cin
-- Output signals: R
--  approx. input signal timings: X: (c11, 0.465385ns)Y: (c11, 0.465385ns)Cin: (c0, 0.000000ns)
--  approx. output signal timings: R: (c11, 1.735385ns)

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntAdder_28_Freq500_uid60 is
    port (clk : in std_logic;
          X : in  std_logic_vector(27 downto 0);
          Y : in  std_logic_vector(27 downto 0);
          Cin : in  std_logic;
          R : out  std_logic_vector(27 downto 0)   );
end entity;

architecture arch of IntAdder_28_Freq500_uid60 is
signal Rtmp :  std_logic_vector(27 downto 0);
   -- timing of Rtmp: (c11, 1.735385ns)
signal Cin_d1, Cin_d2, Cin_d3, Cin_d4, Cin_d5, Cin_d6, Cin_d7, Cin_d8, Cin_d9, Cin_d10, Cin_d11 :  std_logic;
   -- timing of Cin: (c0, 0.000000ns)
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            Cin_d1 <=  Cin;
            Cin_d2 <=  Cin_d1;
            Cin_d3 <=  Cin_d2;
            Cin_d4 <=  Cin_d3;
            Cin_d5 <=  Cin_d4;
            Cin_d6 <=  Cin_d5;
            Cin_d7 <=  Cin_d6;
            Cin_d8 <=  Cin_d7;
            Cin_d9 <=  Cin_d8;
            Cin_d10 <=  Cin_d9;
            Cin_d11 <=  Cin_d10;
         end if;
      end process;
   Rtmp <= X + Y + Cin_d11;
   R <= Rtmp;
end architecture;

--------------------------------------------------------------------------------
--                   FPLogIterative_8_20_0_500_Freq500_uid9
-- VHDL generated for DummyFPGA @ 500MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: F. de Dinechin, C. Klein  (2008-2011)
--------------------------------------------------------------------------------
-- Pipeline depth: 11 cycles
-- Clock period (ns): 2
-- Target frequency (MHz): 500
-- Input signals: X
-- Output signals: R
--  approx. input signal timings: X: (c0, 0.000000ns)
--  approx. output signal timings: R: (c11, 1.735385ns)

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity FPLogIterative_8_20_0_500_Freq500_uid9 is
    port (clk : in std_logic;
          X : in  std_logic_vector(8+20+2 downto 0);
          R : out  std_logic_vector(8+20+2 downto 0)   );
end entity;

architecture arch of FPLogIterative_8_20_0_500_Freq500_uid9 is
   component LZOC_20_Freq500_uid11 is
      port ( clk : in std_logic;
             I : in  std_logic_vector(19 downto 0);
             OZB : in  std_logic;
             O : out  std_logic_vector(4 downto 0)   );
   end component;

   component LeftShifter11_by_max_11_Freq500_uid13 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(10 downto 0);
             S : in  std_logic_vector(3 downto 0);
             R : out  std_logic_vector(21 downto 0)   );
   end component;

   component InvA0Table_Freq500_uid15 is
      port ( X : in  std_logic_vector(7 downto 0);
             Y : out  std_logic_vector(8 downto 0)   );
   end component;

   component IntAdder_24_Freq500_uid19 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(23 downto 0);
             Y : in  std_logic_vector(23 downto 0);
             Cin : in  std_logic;
             R : out  std_logic_vector(23 downto 0)   );
   end component;

   component IntAdder_24_Freq500_uid22 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(23 downto 0);
             Y : in  std_logic_vector(23 downto 0);
             Cin : in  std_logic;
             R : out  std_logic_vector(23 downto 0)   );
   end component;

   component IntAdder_24_Freq500_uid25 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(23 downto 0);
             Y : in  std_logic_vector(23 downto 0);
             Cin : in  std_logic;
             R : out  std_logic_vector(23 downto 0)   );
   end component;

   component LogTable0_Freq500_uid27 is
      port ( X : in  std_logic_vector(7 downto 0);
             Y : out  std_logic_vector(34 downto 0)   );
   end component;

   component LogTable1_Freq500_uid30 is
      port ( X : in  std_logic_vector(5 downto 0);
             Y : out  std_logic_vector(28 downto 0)   );
   end component;

   component IntAdder_35_Freq500_uid34 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(34 downto 0);
             Y : in  std_logic_vector(34 downto 0);
             Cin : in  std_logic;
             R : out  std_logic_vector(34 downto 0)   );
   end component;

   component IntAdder_35_Freq500_uid37 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(34 downto 0);
             Y : in  std_logic_vector(34 downto 0);
             Cin : in  std_logic;
             R : out  std_logic_vector(34 downto 0)   );
   end component;

   component FixRealKCM_Freq500_uid39 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(7 downto 0);
             R : out  std_logic_vector(31 downto 0)   );
   end component;

   component IntAdder_43_Freq500_uid51 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(42 downto 0);
             Y : in  std_logic_vector(42 downto 0);
             Cin : in  std_logic;
             R : out  std_logic_vector(42 downto 0)   );
   end component;

   component Normalizer_Z_43_35_18_Freq500_uid53 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(42 downto 0);
             Count : out  std_logic_vector(4 downto 0);
             R : out  std_logic_vector(34 downto 0)   );
   end component;

   component RightShifter15_by_max_14_Freq500_uid55 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(14 downto 0);
             S : in  std_logic_vector(3 downto 0);
             R : out  std_logic_vector(28 downto 0)   );
   end component;

   component IntAdder_26_Freq500_uid57 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(25 downto 0);
             Y : in  std_logic_vector(25 downto 0);
             Cin : in  std_logic;
             R : out  std_logic_vector(25 downto 0)   );
   end component;

   component IntAdder_28_Freq500_uid60 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(27 downto 0);
             Y : in  std_logic_vector(27 downto 0);
             Cin : in  std_logic;
             R : out  std_logic_vector(27 downto 0)   );
   end component;

signal XExnSgn, XExnSgn_d1, XExnSgn_d2, XExnSgn_d3, XExnSgn_d4, XExnSgn_d5, XExnSgn_d6, XExnSgn_d7, XExnSgn_d8, XExnSgn_d9, XExnSgn_d10, XExnSgn_d11 :  std_logic_vector(2 downto 0);
   -- timing of XExnSgn: (c0, 0.000000ns)
signal FirstBit :  std_logic;
   -- timing of FirstBit: (c0, 0.000000ns)
signal Y0, Y0_d1 :  std_logic_vector(21 downto 0);
   -- timing of Y0: (c0, 0.550000ns)
signal Y0h :  std_logic_vector(19 downto 0);
   -- timing of Y0h: (c0, 0.550000ns)
signal sR, sR_d1, sR_d2, sR_d3, sR_d4, sR_d5, sR_d6, sR_d7, sR_d8, sR_d9, sR_d10, sR_d11 :  std_logic;
   -- timing of sR: (c0, 0.550000ns)
signal absZ0 :  std_logic_vector(10 downto 0);
   -- timing of absZ0: (c0, 1.650000ns)
signal E :  std_logic_vector(7 downto 0);
   -- timing of E: (c0, 1.070000ns)
signal absE :  std_logic_vector(7 downto 0);
   -- timing of absE: (c0, 1.620000ns)
signal EeqZero, EeqZero_d1, EeqZero_d2, EeqZero_d3, EeqZero_d4 :  std_logic;
   -- timing of EeqZero: (c0, 1.620000ns)
signal lzo, lzo_d1, lzo_d2, lzo_d3 :  std_logic_vector(4 downto 0);
   -- timing of lzo: (c3, 0.410000ns)
signal pfinal_s, pfinal_s_d1, pfinal_s_d2, pfinal_s_d3 :  std_logic_vector(4 downto 0);
   -- timing of pfinal_s: (c0, 0.000000ns)
signal shiftval :  std_logic_vector(5 downto 0);
   -- timing of shiftval: (c3, 1.460000ns)
signal shiftvalinL :  std_logic_vector(3 downto 0);
   -- timing of shiftvalinL: (c3, 1.460000ns)
signal shiftvalinR :  std_logic_vector(3 downto 0);
   -- timing of shiftvalinR: (c3, 1.460000ns)
signal doRR, doRR_d1, doRR_d2 :  std_logic;
   -- timing of doRR: (c3, 1.460000ns)
signal small, small_d1, small_d2, small_d3, small_d4, small_d5, small_d6, small_d7 :  std_logic;
   -- timing of small: (c4, 0.210000ns)
signal small_absZ0_normd_full :  std_logic_vector(21 downto 0);
   -- timing of small_absZ0_normd_full: (c4, 1.375385ns)
signal small_absZ0_normd, small_absZ0_normd_d1 :  std_logic_vector(10 downto 0);
   -- timing of small_absZ0_normd: (c4, 1.375385ns)
signal A0 :  std_logic_vector(7 downto 0);
   -- timing of A0: (c0, 0.000000ns)
signal InvA0, InvA0_d1 :  std_logic_vector(8 downto 0);
   -- timing of InvA0: (c0, 0.550000ns)
signal InvA0_copy16 :  std_logic_vector(8 downto 0);
   -- timing of InvA0_copy16: (c0, 0.000000ns)
signal P0 :  std_logic_vector(30 downto 0);
   -- timing of P0: (c1, 0.600000ns)
signal Z1 :  std_logic_vector(22 downto 0);
   -- timing of Z1: (c1, 0.600000ns)
signal A1, A1_d1 :  std_logic_vector(5 downto 0);
   -- timing of A1: (c1, 0.600000ns)
signal B1 :  std_logic_vector(16 downto 0);
   -- timing of B1: (c1, 0.600000ns)
signal ZM1, ZM1_d1 :  std_logic_vector(22 downto 0);
   -- timing of ZM1: (c1, 0.600000ns)
signal P1 :  std_logic_vector(28 downto 0);
   -- timing of P1: (c2, 0.630000ns)
signal Y1 :  std_logic_vector(29 downto 0);
   -- timing of Y1: (c1, 0.600000ns)
signal EiY1 :  std_logic_vector(23 downto 0);
   -- timing of EiY1: (c1, 1.150000ns)
signal addXIter1 :  std_logic_vector(23 downto 0);
   -- timing of addXIter1: (c1, 0.600000ns)
signal EiYPB1 :  std_logic_vector(23 downto 0);
   -- timing of EiYPB1: (c2, 0.590000ns)
signal Pp1 :  std_logic_vector(23 downto 0);
   -- timing of Pp1: (c2, 1.180000ns)
signal Z2 :  std_logic_vector(23 downto 0);
   -- timing of Z2: (c3, 0.620000ns)
signal Zfinal, Zfinal_d1, Zfinal_d2 :  std_logic_vector(23 downto 0);
   -- timing of Zfinal: (c3, 0.620000ns)
signal squarerIn :  std_logic_vector(14 downto 0);
   -- timing of squarerIn: (c5, 0.125385ns)
signal Z2o2_full :  std_logic_vector(29 downto 0);
   -- timing of Z2o2_full: (c5, 0.125385ns)
signal Z2o2_full_dummy :  std_logic_vector(29 downto 0);
   -- timing of Z2o2_full_dummy: (c5, 0.125385ns)
signal Z2o2_normal :  std_logic_vector(11 downto 0);
   -- timing of Z2o2_normal: (c5, 0.125385ns)
signal addFinalLog1pY :  std_logic_vector(23 downto 0);
   -- timing of addFinalLog1pY: (c5, 0.675385ns)
signal Log1p_normal :  std_logic_vector(23 downto 0);
   -- timing of Log1p_normal: (c6, 0.105385ns)
signal L0 :  std_logic_vector(34 downto 0);
   -- timing of L0: (c0, 0.550000ns)
signal L0_copy28 :  std_logic_vector(34 downto 0);
   -- timing of L0_copy28: (c0, 0.000000ns)
signal S1 :  std_logic_vector(34 downto 0);
   -- timing of S1: (c0, 0.550000ns)
signal L1 :  std_logic_vector(28 downto 0);
   -- timing of L1: (c1, 1.200000ns)
signal L1_copy31 :  std_logic_vector(28 downto 0);
   -- timing of L1_copy31: (c1, 0.600000ns)
signal sopX1 :  std_logic_vector(34 downto 0);
   -- timing of sopX1: (c1, 1.200000ns)
signal S2 :  std_logic_vector(34 downto 0);
   -- timing of S2: (c2, 0.750000ns)
signal almostLog :  std_logic_vector(34 downto 0);
   -- timing of almostLog: (c2, 0.750000ns)
signal adderLogF_normalY :  std_logic_vector(34 downto 0);
   -- timing of adderLogF_normalY: (c6, 0.105385ns)
signal LogF_normal :  std_logic_vector(34 downto 0);
   -- timing of LogF_normal: (c6, 1.445385ns)
signal absELog2 :  std_logic_vector(31 downto 0);
   -- timing of absELog2: (c1, 1.680000ns)
signal absELog2_pad :  std_logic_vector(42 downto 0);
   -- timing of absELog2_pad: (c1, 1.680000ns)
signal LogF_normal_pad :  std_logic_vector(42 downto 0);
   -- timing of LogF_normal_pad: (c6, 1.445385ns)
signal lnaddX :  std_logic_vector(42 downto 0);
   -- timing of lnaddX: (c1, 1.680000ns)
signal lnaddY :  std_logic_vector(42 downto 0);
   -- timing of lnaddY: (c6, 1.445385ns)
signal Log_normal :  std_logic_vector(42 downto 0);
   -- timing of Log_normal: (c8, 0.275385ns)
signal Log_normal_normd :  std_logic_vector(34 downto 0);
   -- timing of Log_normal_normd: (c11, 0.465385ns)
signal E_normal :  std_logic_vector(4 downto 0);
   -- timing of E_normal: (c10, 1.715385ns)
signal Z2o2_small_bs :  std_logic_vector(14 downto 0);
   -- timing of Z2o2_small_bs: (c5, 0.125385ns)
signal Z2o2_small_s :  std_logic_vector(28 downto 0);
   -- timing of Z2o2_small_s: (c6, 0.163846ns)
signal Z2o2_small :  std_logic_vector(25 downto 0);
   -- timing of Z2o2_small: (c6, 0.163846ns)
signal Z_small :  std_logic_vector(25 downto 0);
   -- timing of Z_small: (c4, 1.375385ns)
signal Log_smallY :  std_logic_vector(25 downto 0);
   -- timing of Log_smallY: (c6, 0.163846ns)
signal nsRCin :  std_logic;
   -- timing of nsRCin: (c0, 0.550000ns)
signal Log_small :  std_logic_vector(25 downto 0);
   -- timing of Log_small: (c6, 1.413846ns)
signal E0_sub :  std_logic_vector(1 downto 0);
   -- timing of E0_sub: (c6, 1.413846ns)
signal ufl, ufl_d1, ufl_d2, ufl_d3, ufl_d4, ufl_d5, ufl_d6, ufl_d7, ufl_d8, ufl_d9, ufl_d10, ufl_d11 :  std_logic;
   -- timing of ufl: (c0, 0.000000ns)
signal E_small, E_small_d1, E_small_d2, E_small_d3, E_small_d4 :  std_logic_vector(7 downto 0);
   -- timing of E_small: (c6, 1.413846ns)
signal Log_small_normd, Log_small_normd_d1, Log_small_normd_d2, Log_small_normd_d3, Log_small_normd_d4, Log_small_normd_d5 :  std_logic_vector(23 downto 0);
   -- timing of Log_small_normd: (c6, 1.413846ns)
signal E0offset, E0offset_d1, E0offset_d2, E0offset_d3, E0offset_d4, E0offset_d5, E0offset_d6, E0offset_d7, E0offset_d8, E0offset_d9, E0offset_d10 :  std_logic_vector(7 downto 0);
   -- timing of E0offset: (c0, 0.000000ns)
signal ER, ER_d1 :  std_logic_vector(7 downto 0);
   -- timing of ER: (c10, 1.715385ns)
signal Log_g :  std_logic_vector(23 downto 0);
   -- timing of Log_g: (c11, 0.465385ns)
signal round :  std_logic;
   -- timing of round: (c11, 0.465385ns)
signal fraX :  std_logic_vector(27 downto 0);
   -- timing of fraX: (c11, 0.465385ns)
signal fraY :  std_logic_vector(27 downto 0);
   -- timing of fraY: (c11, 0.465385ns)
signal EFR :  std_logic_vector(27 downto 0);
   -- timing of EFR: (c11, 1.735385ns)
signal Rexn :  std_logic_vector(2 downto 0);
   -- timing of Rexn: (c11, 1.015385ns)
constant g: positive := 4;
constant log2wF: positive := 5;
constant pfinal: positive := 11;
constant sfinal: positive := 24;
constant targetprec: positive := 35;
constant wE: positive := 8;
constant wF: positive := 20;
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            XExnSgn_d1 <=  XExnSgn;
            XExnSgn_d2 <=  XExnSgn_d1;
            XExnSgn_d3 <=  XExnSgn_d2;
            XExnSgn_d4 <=  XExnSgn_d3;
            XExnSgn_d5 <=  XExnSgn_d4;
            XExnSgn_d6 <=  XExnSgn_d5;
            XExnSgn_d7 <=  XExnSgn_d6;
            XExnSgn_d8 <=  XExnSgn_d7;
            XExnSgn_d9 <=  XExnSgn_d8;
            XExnSgn_d10 <=  XExnSgn_d9;
            XExnSgn_d11 <=  XExnSgn_d10;
            Y0_d1 <=  Y0;
            sR_d1 <=  sR;
            sR_d2 <=  sR_d1;
            sR_d3 <=  sR_d2;
            sR_d4 <=  sR_d3;
            sR_d5 <=  sR_d4;
            sR_d6 <=  sR_d5;
            sR_d7 <=  sR_d6;
            sR_d8 <=  sR_d7;
            sR_d9 <=  sR_d8;
            sR_d10 <=  sR_d9;
            sR_d11 <=  sR_d10;
            EeqZero_d1 <=  EeqZero;
            EeqZero_d2 <=  EeqZero_d1;
            EeqZero_d3 <=  EeqZero_d2;
            EeqZero_d4 <=  EeqZero_d3;
            lzo_d1 <=  lzo;
            lzo_d2 <=  lzo_d1;
            lzo_d3 <=  lzo_d2;
            pfinal_s_d1 <=  pfinal_s;
            pfinal_s_d2 <=  pfinal_s_d1;
            pfinal_s_d3 <=  pfinal_s_d2;
            doRR_d1 <=  doRR;
            doRR_d2 <=  doRR_d1;
            small_d1 <=  small;
            small_d2 <=  small_d1;
            small_d3 <=  small_d2;
            small_d4 <=  small_d3;
            small_d5 <=  small_d4;
            small_d6 <=  small_d5;
            small_d7 <=  small_d6;
            small_absZ0_normd_d1 <=  small_absZ0_normd;
            InvA0_d1 <=  InvA0;
            A1_d1 <=  A1;
            ZM1_d1 <=  ZM1;
            Zfinal_d1 <=  Zfinal;
            Zfinal_d2 <=  Zfinal_d1;
            ufl_d1 <=  ufl;
            ufl_d2 <=  ufl_d1;
            ufl_d3 <=  ufl_d2;
            ufl_d4 <=  ufl_d3;
            ufl_d5 <=  ufl_d4;
            ufl_d6 <=  ufl_d5;
            ufl_d7 <=  ufl_d6;
            ufl_d8 <=  ufl_d7;
            ufl_d9 <=  ufl_d8;
            ufl_d10 <=  ufl_d9;
            ufl_d11 <=  ufl_d10;
            E_small_d1 <=  E_small;
            E_small_d2 <=  E_small_d1;
            E_small_d3 <=  E_small_d2;
            E_small_d4 <=  E_small_d3;
            Log_small_normd_d1 <=  Log_small_normd;
            Log_small_normd_d2 <=  Log_small_normd_d1;
            Log_small_normd_d3 <=  Log_small_normd_d2;
            Log_small_normd_d4 <=  Log_small_normd_d3;
            Log_small_normd_d5 <=  Log_small_normd_d4;
            E0offset_d1 <=  E0offset;
            E0offset_d2 <=  E0offset_d1;
            E0offset_d3 <=  E0offset_d2;
            E0offset_d4 <=  E0offset_d3;
            E0offset_d5 <=  E0offset_d4;
            E0offset_d6 <=  E0offset_d5;
            E0offset_d7 <=  E0offset_d6;
            E0offset_d8 <=  E0offset_d7;
            E0offset_d9 <=  E0offset_d8;
            E0offset_d10 <=  E0offset_d9;
            ER_d1 <=  ER;
         end if;
      end process;
   XExnSgn <=  X(wE+wF+2 downto wE+wF);
   FirstBit <=  X(wF-1);
   Y0 <= "1" & X(wF-1 downto 0) & "0" when FirstBit = '0' else "01" & X(wF-1 downto 0);
   Y0h <= Y0(wF downto 1);
   -- Sign of the result;
   sR <= '0'   when  (X(wE+wF-1 downto wF) = ('0' & (wE-2 downto 0 => '1')))  -- binade [1..2)
     else not X(wE+wF-1);                -- MSB of exponent
   absZ0 <=   Y0(wF-pfinal+1 downto 0)          when (sR='0') else
             ((wF-pfinal+1 downto 0 => '0') - Y0(wF-pfinal+1 downto 0));
   E <= (X(wE+wF-1 downto wF)) - ("0" & (wE-2 downto 1 => '1') & (not FirstBit));
   absE <= ((wE-1 downto 0 => '0') - E)   when sR = '1' else E;
   EeqZero <= '1' when E=(wE-1 downto 0 => '0') else '0';
   lzoc1: LZOC_20_Freq500_uid11
      port map ( clk  => clk,
                 I => Y0h,
                 OZB => FirstBit,
                 O => lzo);
   pfinal_s <= "01011";
   shiftval <= ('0' & lzo) - ('0' & pfinal_s_d3); 
   shiftvalinL <= shiftval(3 downto 0);
   shiftvalinR <= shiftval(3 downto 0);
   doRR <= shiftval(log2wF); -- sign of the result
   small <= EeqZero_d4 and not(doRR_d1);
   -- The left shifter for the 'small' case
   small_lshift: LeftShifter11_by_max_11_Freq500_uid13
      port map ( clk  => clk,
                 S => shiftvalinL,
                 X => absZ0,
                 R => small_absZ0_normd_full);
   small_absZ0_normd <= small_absZ0_normd_full(10 downto 0); -- get rid of leading zeroes
   ---------------- The range reduction box ---------------
   A0 <= X(19 downto 12);
   -- First inv table
   InvA0Table: InvA0Table_Freq500_uid15
      port map ( X => A0,
                 Y => InvA0_copy16);
   InvA0 <= InvA0_copy16; -- output copy to hold a pipeline register if needed
   P0 <= InvA0_d1 * Y0_d1;

   Z1 <= P0(22 downto 0);

   A1 <= Z1(22 downto 17);
   B1 <= Z1(16 downto 0);
   ZM1 <= Z1;
   P1 <= A1_d1*ZM1_d1;
   Y1 <= "1" & (5 downto 0 => '0') & Z1;
   EiY1 <= Y1(29 downto 6)  when A1(5) = '1'
     else  "0" & Y1(29 downto 7);
   addXIter1 <= "0" & B1 & (5 downto 0 => '0');
   addIter1_1: IntAdder_24_Freq500_uid19
      port map ( clk  => clk,
                 Cin => '0',
                 X => addXIter1,
                 Y => EiY1,
                 R => EiYPB1);
   Pp1 <= (0 downto 0 => '1') & not(P1(28 downto 6));
   addIter2_1: IntAdder_24_Freq500_uid22
      port map ( clk  => clk,
                 Cin => '1',
                 X => EiYPB1,
                 Y => Pp1,
                 R => Z2);
   Zfinal <= Z2;
   squarerIn <= Zfinal_d2(sfinal-1 downto sfinal-15) when doRR_d2='1'
                    else (small_absZ0_normd_d1 & (3 downto 0 => '0'));  
   Z2o2_full <= squarerIn*squarerIn;
   Z2o2_full_dummy <= Z2o2_full;
   Z2o2_normal <= Z2o2_full_dummy (29  downto 18);
   addFinalLog1pY <= (pfinal downto 0  => '1') & not(Z2o2_normal);
   addFinalLog1p_normalAdder: IntAdder_24_Freq500_uid25
      port map ( clk  => clk,
                 Cin => '1',
                 X => Zfinal,
                 Y => addFinalLog1pY,
                 R => Log1p_normal);

   -- Now the log tables, as late as possible
   LogTable0: LogTable0_Freq500_uid27
      port map ( X => A0,
                 Y => L0_copy28);
   L0 <= L0_copy28; -- output copy to hold a pipeline register if needed
   S1 <= L0;
   LogTable1: LogTable1_Freq500_uid30
      port map ( X => A1,
                 Y => L1_copy31);
   L1 <= L1_copy31; -- output copy to hold a pipeline register if needed
   sopX1 <= ((34 downto 29 => '0') & L1);
   adderS1: IntAdder_35_Freq500_uid34
      port map ( clk  => clk,
                 Cin => '0',
                 X => S1,
                 Y => sopX1,
                 R => S2);
   almostLog <= S2;
   adderLogF_normalY <= ((targetprec-1 downto sfinal => '0') & Log1p_normal);
   adderLogF_normal: IntAdder_35_Freq500_uid37
      port map ( clk  => clk,
                 Cin => '0',
                 X => almostLog,
                 Y => adderLogF_normalY,
                 R => LogF_normal);
   MulLog2: FixRealKCM_Freq500_uid39
      port map ( clk  => clk,
                 X => absE,
                 R => absELog2);
   absELog2_pad <=   absELog2 & (targetprec-wF-g-1 downto 0 => '0');       
   LogF_normal_pad <= (wE-1  downto 0 => LogF_normal(targetprec-1))  & LogF_normal;
   lnaddX <= absELog2_pad;
   lnaddY <= LogF_normal_pad when sR_d6='0' else not(LogF_normal_pad); 
   lnadder: IntAdder_43_Freq500_uid51
      port map ( clk  => clk,
                 Cin => sR,
                 X => lnaddX,
                 Y => lnaddY,
                 R => Log_normal);
   final_norm: Normalizer_Z_43_35_18_Freq500_uid53
      port map ( clk  => clk,
                 X => Log_normal,
                 Count => E_normal,
                 R => Log_normal_normd);
   Z2o2_small_bs <= Z2o2_full_dummy(29 downto 15);
   ao_rshift: RightShifter15_by_max_14_Freq500_uid55
      port map ( clk  => clk,
                 S => shiftvalinR,
                 X => Z2o2_small_bs,
                 R => Z2o2_small_s);
     -- send the MSB to position pfinal
   Z2o2_small <=  (pfinal-1 downto 0  => '0') & Z2o2_small_s(28 downto 14);
   -- mantissa will be either Y0-z^2/2  or  -Y0+z^2/2,  depending on sR  
   Z_small <= small_absZ0_normd & (14 downto 0 => '0');
   Log_smallY <= Z2o2_small when sR_d6='1' else not(Z2o2_small);
   nsRCin <= not ( sR );
   log_small_adder: IntAdder_26_Freq500_uid57
      port map ( clk  => clk,
                 Cin => nsRCin,
                 X => Z_small,
                 Y => Log_smallY,
                 R => Log_small);
   -- Possibly subtract 1 or 2 to the exponent, depending on the LZC of Log_small
   E0_sub <=   "11" when Log_small(wF+g+1) = '1'
          else "10" when Log_small(wF+g+1 downto wF+g) = "01"
          else "01" ;
   -- The smallest log will be log(1+2^{-wF}) \approx 2^{-wF}  = 2^-20
   -- The smallest representable number is 2^{1-2^(wE-1)} = 2^-127
   -- No underflow possible
   ufl <= '0';
   E_small <=  ("0" & (wE-2 downto 2 => '1') & E0_sub)  -  ((wE-1 downto 5 => '0') & lzo_d3) ;
   Log_small_normd <= Log_small(wF+g+1 downto 2) when Log_small(wF+g+1)='1'
           else Log_small(wF+g downto 1)  when Log_small(wF+g)='1'  -- remove the first zero
           else Log_small(wF+g-1 downto 0)  ; -- remove two zeroes (extremely rare, 001000000 only)
   E0offset <= "10000110"; -- E0 + wE 
   ER <= E_small_d4(7 downto 0) when small_d6='1'
      else E0offset_d10 - ((7 downto 5 => '0') & E_normal);
   Log_g <=  Log_small_normd_d5(wF+g-2 downto 0) & "0" when small_d7='1'           -- remove implicit 1
      else Log_normal_normd(targetprec-2 downto targetprec-wF-g-1 );  -- remove implicit 1
   round <= Log_g(g-1) ; -- sticky is always 1 for a transcendental function 
   -- if round leads to a change of binade, the carry propagation magically updates both mantissa and exponent
   fraX <= (ER_d1 & Log_g(wF+g-1 downto g)) ; 
   fraY <= ((wE+wF-1 downto 1 => '0') & round); 
   finalRoundAdder: IntAdder_28_Freq500_uid60
      port map ( clk  => clk,
                 Cin => '0',
                 X => fraX,
                 Y => fraY,
                 R => EFR);
   Rexn <= "110" when ((XExnSgn_d11(2) and (XExnSgn_d11(1) or XExnSgn_d11(0))) or (XExnSgn_d11(1) and XExnSgn_d11(0))) = '1' else
                              "101" when XExnSgn_d11(2 downto 1) = "00"  else
                              "100" when XExnSgn_d11(2 downto 1) = "10"  else
                              "00" & sR_d11 when (((Log_normal_normd(targetprec-1)='0') and (small_d7='0')) or ( (Log_small_normd_d5 (wF+g-1)='0') and (small_d7='1'))) or (ufl_d11 = '1' and small_d7='1') else
                               "01" & sR_d11;
   R<=  Rexn & EFR;
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplier_21x11_24_Freq500_uid65
-- VHDL generated for DummyFPGA @ 500MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Martin Kumm, Florent de Dinechin, Andreas Böttcher, Kinga Illyes, Bogdan Popa, Bogdan Pasca, 2012-
--------------------------------------------------------------------------------
-- Pipeline depth: 11 cycles
-- Clock period (ns): 2
-- Target frequency (MHz): 500
-- Input signals: X Y
-- Output signals: R
--  approx. input signal timings: X: (c11, 1.735385ns)Y: (c0, 0.000000ns)
--  approx. output signal timings: R: (c11, 1.735385ns)

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity IntMultiplier_21x11_24_Freq500_uid65 is
    port (clk : in std_logic;
          X : in  std_logic_vector(20 downto 0);
          Y : in  std_logic_vector(10 downto 0);
          R : out  std_logic_vector(23 downto 0)   );
end entity;

architecture arch of IntMultiplier_21x11_24_Freq500_uid65 is
signal XX_m66 :  std_logic_vector(20 downto 0);
   -- timing of XX_m66: (c11, 1.735385ns)
signal YY_m66 :  std_logic_vector(10 downto 0);
   -- timing of YY_m66: (c0, 0.000000ns)
signal XX :  unsigned(-1+21 downto 0);
   -- timing of XX: (c11, 1.735385ns)
signal YY, YY_d1, YY_d2, YY_d3, YY_d4, YY_d5, YY_d6, YY_d7, YY_d8, YY_d9, YY_d10, YY_d11 :  unsigned(-1+11 downto 0);
   -- timing of YY: (c0, 0.000000ns)
signal RR :  unsigned(-1+32 downto 0);
   -- timing of RR: (c11, 1.735385ns)
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            YY_d1 <=  YY;
            YY_d2 <=  YY_d1;
            YY_d3 <=  YY_d2;
            YY_d4 <=  YY_d3;
            YY_d5 <=  YY_d4;
            YY_d6 <=  YY_d5;
            YY_d7 <=  YY_d6;
            YY_d8 <=  YY_d7;
            YY_d9 <=  YY_d8;
            YY_d10 <=  YY_d9;
            YY_d11 <=  YY_d10;
         end if;
      end process;
   XX_m66 <= X ;
   YY_m66 <= Y ;
   XX <= unsigned(X);
   YY <= unsigned(Y);
   RR <= XX*YY_d11;
   R <= std_logic_vector(RR(31 downto 8));
end architecture;

--------------------------------------------------------------------------------
--                         IntAdder_31_Freq500_uid69
-- VHDL generated for DummyFPGA @ 500MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin (2008-2016)
--------------------------------------------------------------------------------
-- Pipeline depth: 13 cycles
-- Clock period (ns): 2
-- Target frequency (MHz): 500
-- Input signals: X Y Cin
-- Output signals: R
--  approx. input signal timings: X: (c13, 0.315385ns)Y: (c0, 0.000000ns)Cin: (c0, 0.000000ns)
--  approx. output signal timings: R: (c13, 1.615385ns)

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntAdder_31_Freq500_uid69 is
    port (clk : in std_logic;
          X : in  std_logic_vector(30 downto 0);
          Y : in  std_logic_vector(30 downto 0);
          Cin : in  std_logic;
          R : out  std_logic_vector(30 downto 0)   );
end entity;

architecture arch of IntAdder_31_Freq500_uid69 is
signal Rtmp :  std_logic_vector(30 downto 0);
   -- timing of Rtmp: (c13, 1.615385ns)
signal Y_d1, Y_d2, Y_d3, Y_d4, Y_d5, Y_d6, Y_d7, Y_d8, Y_d9, Y_d10, Y_d11, Y_d12, Y_d13 :  std_logic_vector(30 downto 0);
   -- timing of Y: (c0, 0.000000ns)
signal Cin_d1, Cin_d2, Cin_d3, Cin_d4, Cin_d5, Cin_d6, Cin_d7, Cin_d8, Cin_d9, Cin_d10, Cin_d11, Cin_d12, Cin_d13 :  std_logic;
   -- timing of Cin: (c0, 0.000000ns)
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            Y_d1 <=  Y;
            Y_d2 <=  Y_d1;
            Y_d3 <=  Y_d2;
            Y_d4 <=  Y_d3;
            Y_d5 <=  Y_d4;
            Y_d6 <=  Y_d5;
            Y_d7 <=  Y_d6;
            Y_d8 <=  Y_d7;
            Y_d9 <=  Y_d8;
            Y_d10 <=  Y_d9;
            Y_d11 <=  Y_d10;
            Y_d12 <=  Y_d11;
            Y_d13 <=  Y_d12;
            Cin_d1 <=  Cin;
            Cin_d2 <=  Cin_d1;
            Cin_d3 <=  Cin_d2;
            Cin_d4 <=  Cin_d3;
            Cin_d5 <=  Cin_d4;
            Cin_d6 <=  Cin_d5;
            Cin_d7 <=  Cin_d6;
            Cin_d8 <=  Cin_d7;
            Cin_d9 <=  Cin_d8;
            Cin_d10 <=  Cin_d9;
            Cin_d11 <=  Cin_d10;
            Cin_d12 <=  Cin_d11;
            Cin_d13 <=  Cin_d12;
         end if;
      end process;
   Rtmp <= X + Y_d13 + Cin_d13;
   R <= Rtmp;
end architecture;

--------------------------------------------------------------------------------
--                      FPMult_8_20_uid62_Freq500_uid63
-- VHDL generated for DummyFPGA @ 500MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin 2008-2021
--------------------------------------------------------------------------------
-- Pipeline depth: 13 cycles
-- Clock period (ns): 2
-- Target frequency (MHz): 500
-- Input signals: X Y
-- Output signals: R
--  approx. input signal timings: X: (c11, 1.735385ns)Y: (c0, 0.000000ns)
--  approx. output signal timings: R: (c13, 1.615385ns)

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity FPMult_8_20_uid62_Freq500_uid63 is
    port (clk : in std_logic;
          X : in  std_logic_vector(8+20+2 downto 0);
          Y : in  std_logic_vector(8+10+2 downto 0);
          R : out  std_logic_vector(8+21+2 downto 0)   );
end entity;

architecture arch of FPMult_8_20_uid62_Freq500_uid63 is
   component IntMultiplier_21x11_24_Freq500_uid65 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(20 downto 0);
             Y : in  std_logic_vector(10 downto 0);
             R : out  std_logic_vector(23 downto 0)   );
   end component;

   component IntAdder_31_Freq500_uid69 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(30 downto 0);
             Y : in  std_logic_vector(30 downto 0);
             Cin : in  std_logic;
             R : out  std_logic_vector(30 downto 0)   );
   end component;

signal sign, sign_d1, sign_d2 :  std_logic;
   -- timing of sign: (c11, 1.785385ns)
signal expX, expX_d1 :  std_logic_vector(7 downto 0);
   -- timing of expX: (c11, 1.735385ns)
signal expY, expY_d1, expY_d2, expY_d3, expY_d4, expY_d5, expY_d6, expY_d7, expY_d8, expY_d9, expY_d10, expY_d11, expY_d12 :  std_logic_vector(7 downto 0);
   -- timing of expY: (c0, 0.000000ns)
signal expSumPreSub, expSumPreSub_d1 :  std_logic_vector(9 downto 0);
   -- timing of expSumPreSub: (c12, 1.025385ns)
signal bias, bias_d1, bias_d2, bias_d3, bias_d4, bias_d5, bias_d6, bias_d7, bias_d8, bias_d9, bias_d10, bias_d11, bias_d12, bias_d13 :  std_logic_vector(9 downto 0);
   -- timing of bias: (c0, 0.000000ns)
signal expSum :  std_logic_vector(9 downto 0);
   -- timing of expSum: (c13, 0.315385ns)
signal sigX :  std_logic_vector(20 downto 0);
   -- timing of sigX: (c11, 1.735385ns)
signal sigY :  std_logic_vector(10 downto 0);
   -- timing of sigY: (c0, 0.000000ns)
signal sigProd, sigProd_d1 :  std_logic_vector(23 downto 0);
   -- timing of sigProd: (c11, 1.735385ns)
signal excSel :  std_logic_vector(3 downto 0);
   -- timing of excSel: (c11, 1.735385ns)
signal exc, exc_d1, exc_d2 :  std_logic_vector(1 downto 0);
   -- timing of exc: (c11, 1.785385ns)
signal norm, norm_d1, norm_d2 :  std_logic;
   -- timing of norm: (c11, 1.735385ns)
signal expPostNorm :  std_logic_vector(9 downto 0);
   -- timing of expPostNorm: (c13, 0.315385ns)
signal sigProdExt, sigProdExt_d1 :  std_logic_vector(23 downto 0);
   -- timing of sigProdExt: (c12, 0.485385ns)
signal expSig :  std_logic_vector(30 downto 0);
   -- timing of expSig: (c13, 0.315385ns)
signal round :  std_logic;
   -- timing of round: (c0, 0.000000ns)
signal expSigPostRound :  std_logic_vector(30 downto 0);
   -- timing of expSigPostRound: (c13, 1.615385ns)
signal excPostNorm :  std_logic_vector(1 downto 0);
   -- timing of excPostNorm: (c13, 1.615385ns)
signal finalExc :  std_logic_vector(1 downto 0);
   -- timing of finalExc: (c13, 1.615385ns)
signal Y_d1, Y_d2, Y_d3, Y_d4, Y_d5, Y_d6, Y_d7, Y_d8, Y_d9, Y_d10, Y_d11 :  std_logic_vector(8+10+2 downto 0);
   -- timing of Y: (c0, 0.000000ns)
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            sign_d1 <=  sign;
            sign_d2 <=  sign_d1;
            expX_d1 <=  expX;
            expY_d1 <=  expY;
            expY_d2 <=  expY_d1;
            expY_d3 <=  expY_d2;
            expY_d4 <=  expY_d3;
            expY_d5 <=  expY_d4;
            expY_d6 <=  expY_d5;
            expY_d7 <=  expY_d6;
            expY_d8 <=  expY_d7;
            expY_d9 <=  expY_d8;
            expY_d10 <=  expY_d9;
            expY_d11 <=  expY_d10;
            expY_d12 <=  expY_d11;
            expSumPreSub_d1 <=  expSumPreSub;
            bias_d1 <=  bias;
            bias_d2 <=  bias_d1;
            bias_d3 <=  bias_d2;
            bias_d4 <=  bias_d3;
            bias_d5 <=  bias_d4;
            bias_d6 <=  bias_d5;
            bias_d7 <=  bias_d6;
            bias_d8 <=  bias_d7;
            bias_d9 <=  bias_d8;
            bias_d10 <=  bias_d9;
            bias_d11 <=  bias_d10;
            bias_d12 <=  bias_d11;
            bias_d13 <=  bias_d12;
            sigProd_d1 <=  sigProd;
            exc_d1 <=  exc;
            exc_d2 <=  exc_d1;
            norm_d1 <=  norm;
            norm_d2 <=  norm_d1;
            sigProdExt_d1 <=  sigProdExt;
            Y_d1 <=  Y;
            Y_d2 <=  Y_d1;
            Y_d3 <=  Y_d2;
            Y_d4 <=  Y_d3;
            Y_d5 <=  Y_d4;
            Y_d6 <=  Y_d5;
            Y_d7 <=  Y_d6;
            Y_d8 <=  Y_d7;
            Y_d9 <=  Y_d8;
            Y_d10 <=  Y_d9;
            Y_d11 <=  Y_d10;
         end if;
      end process;
   sign <= X(28) xor Y_d11(18);
   expX <= X(27 downto 20);
   expY <= Y(17 downto 10);
   expSumPreSub <= ("00" & expX_d1) + ("00" & expY_d12);
   bias <= CONV_STD_LOGIC_VECTOR(127,10);
   expSum <= expSumPreSub_d1 - bias_d13;
   sigX <= "1" & X(19 downto 0);
   sigY <= "1" & Y(9 downto 0);
   SignificandMultiplication: IntMultiplier_21x11_24_Freq500_uid65
      port map ( clk  => clk,
                 X => sigX,
                 Y => sigY,
                 R => sigProd);
   excSel <= X(30 downto 29) & Y_d11(20 downto 19);
   with excSel  select  
   exc <= "00" when  "0000" | "0001" | "0100", 
          "01" when "0101",
          "10" when "0110" | "1001" | "1010" ,
          "11" when others;
   norm <= sigProd(23);
   -- exponent update
   expPostNorm <= expSum + ("000000000" & norm_d2);
   -- significand normalization shift
   sigProdExt <= sigProd_d1(22 downto 0) & "0" when norm_d1='1' else
                         sigProd_d1(21 downto 0) & "00";
   expSig <= expPostNorm & sigProdExt_d1(23 downto 3);
   round <= '1' ;
   RoundingAdder: IntAdder_31_Freq500_uid69
      port map ( clk  => clk,
                 Cin => round,
                 X => expSig,
                 Y => "0000000000000000000000000000000",
                 R => expSigPostRound);
   with expSigPostRound(30 downto 29)  select 
   excPostNorm <=  "01"  when  "00",
                               "10"             when "01", 
                               "00"             when "11"|"10",
                               "11"             when others;
   with exc_d2  select  
   finalExc <= exc_d2 when  "11"|"10"|"00",
                       excPostNorm when others; 
   R <= finalExc & sign_d2 & expSigPostRound(28 downto 0);
end architecture;

--------------------------------------------------------------------------------
--                   LeftShifter22_by_max_19_Freq500_uid73
-- VHDL generated for DummyFPGA @ 500MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca (2008-2011), Florent de Dinechin (2008-2019)
--------------------------------------------------------------------------------
-- Pipeline depth: 2 cycles
-- Clock period (ns): 2
-- Target frequency (MHz): 500
-- Input signals: X S
-- Output signals: R
--  approx. input signal timings: X: (c13, 1.615385ns)S: (c14, 0.905385ns)
--  approx. output signal timings: R: (c15, 1.159231ns)

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity LeftShifter22_by_max_19_Freq500_uid73 is
    port (clk : in std_logic;
          X : in  std_logic_vector(21 downto 0);
          S : in  std_logic_vector(4 downto 0);
          R : out  std_logic_vector(40 downto 0)   );
end entity;

architecture arch of LeftShifter22_by_max_19_Freq500_uid73 is
signal ps, ps_d1 :  std_logic_vector(4 downto 0);
   -- timing of ps: (c14, 0.905385ns)
signal level0, level0_d1 :  std_logic_vector(21 downto 0);
   -- timing of level0: (c13, 1.615385ns)
signal level1, level1_d1 :  std_logic_vector(22 downto 0);
   -- timing of level1: (c14, 0.905385ns)
signal level2 :  std_logic_vector(24 downto 0);
   -- timing of level2: (c15, 0.040000ns)
signal level3 :  std_logic_vector(28 downto 0);
   -- timing of level3: (c15, 0.040000ns)
signal level4 :  std_logic_vector(36 downto 0);
   -- timing of level4: (c15, 1.159231ns)
signal level5 :  std_logic_vector(52 downto 0);
   -- timing of level5: (c15, 1.159231ns)
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            ps_d1 <=  ps;
            level0_d1 <=  level0;
            level1_d1 <=  level1;
         end if;
      end process;
   ps<= S;
   level0<= X;
   level1<= level0_d1 & (0 downto 0 => '0') when ps(0)= '1' else     (0 downto 0 => '0') & level0_d1;
   level2<= level1_d1 & (1 downto 0 => '0') when ps_d1(1)= '1' else     (1 downto 0 => '0') & level1_d1;
   level3<= level2 & (3 downto 0 => '0') when ps_d1(2)= '1' else     (3 downto 0 => '0') & level2;
   level4<= level3 & (7 downto 0 => '0') when ps_d1(3)= '1' else     (7 downto 0 => '0') & level3;
   level5<= level4 & (15 downto 0 => '0') when ps_d1(4)= '1' else     (15 downto 0 => '0') & level4;
   R <= level5(40 downto 0);
end architecture;

--------------------------------------------------------------------------------
--                         IntAdder_12_Freq500_uid87
-- VHDL generated for DummyFPGA @ 500MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin (2008-2016)
--------------------------------------------------------------------------------
-- Pipeline depth: 16 cycles
-- Clock period (ns): 2
-- Target frequency (MHz): 500
-- Input signals: X Y Cin
-- Output signals: R
--  approx. input signal timings: X: (c15, 1.709231ns)Y: (c15, 1.709231ns)Cin: (c0, 0.000000ns)
--  approx. output signal timings: R: (c16, 1.019231ns)

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntAdder_12_Freq500_uid87 is
    port (clk : in std_logic;
          X : in  std_logic_vector(11 downto 0);
          Y : in  std_logic_vector(11 downto 0);
          Cin : in  std_logic;
          R : out  std_logic_vector(11 downto 0)   );
end entity;

architecture arch of IntAdder_12_Freq500_uid87 is
signal Rtmp :  std_logic_vector(11 downto 0);
   -- timing of Rtmp: (c16, 1.019231ns)
signal X_d1 :  std_logic_vector(11 downto 0);
   -- timing of X: (c15, 1.709231ns)
signal Y_d1 :  std_logic_vector(11 downto 0);
   -- timing of Y: (c15, 1.709231ns)
signal Cin_d1, Cin_d2, Cin_d3, Cin_d4, Cin_d5, Cin_d6, Cin_d7, Cin_d8, Cin_d9, Cin_d10, Cin_d11, Cin_d12, Cin_d13, Cin_d14, Cin_d15, Cin_d16 :  std_logic;
   -- timing of Cin: (c0, 0.000000ns)
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            X_d1 <=  X;
            Y_d1 <=  Y;
            Cin_d1 <=  Cin;
            Cin_d2 <=  Cin_d1;
            Cin_d3 <=  Cin_d2;
            Cin_d4 <=  Cin_d3;
            Cin_d5 <=  Cin_d4;
            Cin_d6 <=  Cin_d5;
            Cin_d7 <=  Cin_d6;
            Cin_d8 <=  Cin_d7;
            Cin_d9 <=  Cin_d8;
            Cin_d10 <=  Cin_d9;
            Cin_d11 <=  Cin_d10;
            Cin_d12 <=  Cin_d11;
            Cin_d13 <=  Cin_d12;
            Cin_d14 <=  Cin_d13;
            Cin_d15 <=  Cin_d14;
            Cin_d16 <=  Cin_d15;
         end if;
      end process;
   Rtmp <= X_d1 + Y_d1 + Cin_d16;
   R <= Rtmp;
end architecture;

--------------------------------------------------------------------------------
--                          FixRealKCM_Freq500_uid77
-- VHDL generated for DummyFPGA @ 500MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin (2007-2016)
--------------------------------------------------------------------------------
-- Pipeline depth: 1 cycles
-- Clock period (ns): 2
-- Target frequency (MHz): 500
-- Input signals: X
-- Output signals: R
--  approx. input signal timings: X: (c15, 1.159231ns)
--  approx. output signal timings: R: (c16, 1.019231ns)

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity FixRealKCM_Freq500_uid77 is
    port (clk : in std_logic;
          X : in  std_logic_vector(9 downto 0);
          R : out  std_logic_vector(7 downto 0)   );
end entity;

architecture arch of FixRealKCM_Freq500_uid77 is
   component FixRealKCM_Freq500_uid77_T0_Freq500_uid80 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(11 downto 0)   );
   end component;

   component FixRealKCM_Freq500_uid77_T1_Freq500_uid83 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(6 downto 0)   );
   end component;

   component IntAdder_12_Freq500_uid87 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(11 downto 0);
             Y : in  std_logic_vector(11 downto 0);
             Cin : in  std_logic;
             R : out  std_logic_vector(11 downto 0)   );
   end component;

signal FixRealKCM_Freq500_uid77_A0 :  std_logic_vector(4 downto 0);
   -- timing of FixRealKCM_Freq500_uid77_A0: (c15, 1.159231ns)
signal FixRealKCM_Freq500_uid77_T0 :  std_logic_vector(11 downto 0);
   -- timing of FixRealKCM_Freq500_uid77_T0: (c15, 1.709231ns)
signal FixRealKCM_Freq500_uid77_T0_copy81 :  std_logic_vector(11 downto 0);
   -- timing of FixRealKCM_Freq500_uid77_T0_copy81: (c15, 1.159231ns)
signal bh78_w0_0 :  std_logic;
   -- timing of bh78_w0_0: (c15, 1.709231ns)
signal bh78_w1_0 :  std_logic;
   -- timing of bh78_w1_0: (c15, 1.709231ns)
signal bh78_w2_0 :  std_logic;
   -- timing of bh78_w2_0: (c15, 1.709231ns)
signal bh78_w3_0 :  std_logic;
   -- timing of bh78_w3_0: (c15, 1.709231ns)
signal bh78_w4_0 :  std_logic;
   -- timing of bh78_w4_0: (c15, 1.709231ns)
signal bh78_w5_0 :  std_logic;
   -- timing of bh78_w5_0: (c15, 1.709231ns)
signal bh78_w6_0 :  std_logic;
   -- timing of bh78_w6_0: (c15, 1.709231ns)
signal bh78_w7_0 :  std_logic;
   -- timing of bh78_w7_0: (c15, 1.709231ns)
signal bh78_w8_0 :  std_logic;
   -- timing of bh78_w8_0: (c15, 1.709231ns)
signal bh78_w9_0 :  std_logic;
   -- timing of bh78_w9_0: (c15, 1.709231ns)
signal bh78_w10_0 :  std_logic;
   -- timing of bh78_w10_0: (c15, 1.709231ns)
signal bh78_w11_0 :  std_logic;
   -- timing of bh78_w11_0: (c15, 1.709231ns)
signal FixRealKCM_Freq500_uid77_A1 :  std_logic_vector(4 downto 0);
   -- timing of FixRealKCM_Freq500_uid77_A1: (c15, 1.159231ns)
signal FixRealKCM_Freq500_uid77_T1 :  std_logic_vector(6 downto 0);
   -- timing of FixRealKCM_Freq500_uid77_T1: (c15, 1.709231ns)
signal FixRealKCM_Freq500_uid77_T1_copy84 :  std_logic_vector(6 downto 0);
   -- timing of FixRealKCM_Freq500_uid77_T1_copy84: (c15, 1.159231ns)
signal bh78_w0_1 :  std_logic;
   -- timing of bh78_w0_1: (c15, 1.709231ns)
signal bh78_w1_1 :  std_logic;
   -- timing of bh78_w1_1: (c15, 1.709231ns)
signal bh78_w2_1 :  std_logic;
   -- timing of bh78_w2_1: (c15, 1.709231ns)
signal bh78_w3_1 :  std_logic;
   -- timing of bh78_w3_1: (c15, 1.709231ns)
signal bh78_w4_1 :  std_logic;
   -- timing of bh78_w4_1: (c15, 1.709231ns)
signal bh78_w5_1 :  std_logic;
   -- timing of bh78_w5_1: (c15, 1.709231ns)
signal bh78_w6_1 :  std_logic;
   -- timing of bh78_w6_1: (c15, 1.709231ns)
signal bitheapFinalAdd_bh78_In0 :  std_logic_vector(11 downto 0);
   -- timing of bitheapFinalAdd_bh78_In0: (c15, 1.709231ns)
signal bitheapFinalAdd_bh78_In1 :  std_logic_vector(11 downto 0);
   -- timing of bitheapFinalAdd_bh78_In1: (c15, 1.709231ns)
signal bitheapFinalAdd_bh78_Cin :  std_logic;
   -- timing of bitheapFinalAdd_bh78_Cin: (c0, 0.000000ns)
signal bitheapFinalAdd_bh78_Out :  std_logic_vector(11 downto 0);
   -- timing of bitheapFinalAdd_bh78_Out: (c16, 1.019231ns)
signal bitheapResult_bh78 :  std_logic_vector(11 downto 0);
   -- timing of bitheapResult_bh78: (c16, 1.019231ns)
signal OutRes :  std_logic_vector(11 downto 0);
   -- timing of OutRes: (c16, 1.019231ns)
begin
-- This operator multiplies by 1/log(2)
   FixRealKCM_Freq500_uid77_A0 <= X(9 downto 5);-- input address  m=6  l=2
   FixRealKCM_Freq500_uid77_Table0: FixRealKCM_Freq500_uid77_T0_Freq500_uid80
      port map ( X => FixRealKCM_Freq500_uid77_A0,
                 Y => FixRealKCM_Freq500_uid77_T0_copy81);
   FixRealKCM_Freq500_uid77_T0 <= FixRealKCM_Freq500_uid77_T0_copy81; -- output copy to hold a pipeline register if needed
   bh78_w0_0 <= FixRealKCM_Freq500_uid77_T0(0);
   bh78_w1_0 <= FixRealKCM_Freq500_uid77_T0(1);
   bh78_w2_0 <= FixRealKCM_Freq500_uid77_T0(2);
   bh78_w3_0 <= FixRealKCM_Freq500_uid77_T0(3);
   bh78_w4_0 <= FixRealKCM_Freq500_uid77_T0(4);
   bh78_w5_0 <= FixRealKCM_Freq500_uid77_T0(5);
   bh78_w6_0 <= FixRealKCM_Freq500_uid77_T0(6);
   bh78_w7_0 <= FixRealKCM_Freq500_uid77_T0(7);
   bh78_w8_0 <= FixRealKCM_Freq500_uid77_T0(8);
   bh78_w9_0 <= FixRealKCM_Freq500_uid77_T0(9);
   bh78_w10_0 <= FixRealKCM_Freq500_uid77_T0(10);
   bh78_w11_0 <= FixRealKCM_Freq500_uid77_T0(11);
   FixRealKCM_Freq500_uid77_A1 <= X(4 downto 0);-- input address  m=1  l=-3
   FixRealKCM_Freq500_uid77_Table1: FixRealKCM_Freq500_uid77_T1_Freq500_uid83
      port map ( X => FixRealKCM_Freq500_uid77_A1,
                 Y => FixRealKCM_Freq500_uid77_T1_copy84);
   FixRealKCM_Freq500_uid77_T1 <= FixRealKCM_Freq500_uid77_T1_copy84; -- output copy to hold a pipeline register if needed
   bh78_w0_1 <= FixRealKCM_Freq500_uid77_T1(0);
   bh78_w1_1 <= FixRealKCM_Freq500_uid77_T1(1);
   bh78_w2_1 <= FixRealKCM_Freq500_uid77_T1(2);
   bh78_w3_1 <= FixRealKCM_Freq500_uid77_T1(3);
   bh78_w4_1 <= FixRealKCM_Freq500_uid77_T1(4);
   bh78_w5_1 <= FixRealKCM_Freq500_uid77_T1(5);
   bh78_w6_1 <= FixRealKCM_Freq500_uid77_T1(6);

   -- Adding the constant bits 
      -- All the constant bits are zero, nothing to add


   bitheapFinalAdd_bh78_In0 <= "" & bh78_w11_0 & bh78_w10_0 & bh78_w9_0 & bh78_w8_0 & bh78_w7_0 & bh78_w6_0 & bh78_w5_0 & bh78_w4_0 & bh78_w3_0 & bh78_w2_0 & bh78_w1_0 & bh78_w0_0;
   bitheapFinalAdd_bh78_In1 <= "0" & "0" & "0" & "0" & "0" & bh78_w6_1 & bh78_w5_1 & bh78_w4_1 & bh78_w3_1 & bh78_w2_1 & bh78_w1_1 & bh78_w0_1;
   bitheapFinalAdd_bh78_Cin <= '0';

   bitheapFinalAdd_bh78: IntAdder_12_Freq500_uid87
      port map ( clk  => clk,
                 Cin => bitheapFinalAdd_bh78_Cin,
                 X => bitheapFinalAdd_bh78_In0,
                 Y => bitheapFinalAdd_bh78_In1,
                 R => bitheapFinalAdd_bh78_Out);
   bitheapResult_bh78 <= bitheapFinalAdd_bh78_Out(11 downto 0);
   OutRes <= bitheapResult_bh78(11 downto 0);
   R <= OutRes(11 downto 4);
end architecture;

--------------------------------------------------------------------------------
--                         IntAdder_21_Freq500_uid99
-- VHDL generated for DummyFPGA @ 500MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin (2008-2016)
--------------------------------------------------------------------------------
-- Pipeline depth: 17 cycles
-- Clock period (ns): 2
-- Target frequency (MHz): 500
-- Input signals: X Y Cin
-- Output signals: R
--  approx. input signal timings: X: (c16, 1.569231ns)Y: (c16, 1.569231ns)Cin: (c0, 0.000000ns)
--  approx. output signal timings: R: (c17, 0.969231ns)

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntAdder_21_Freq500_uid99 is
    port (clk : in std_logic;
          X : in  std_logic_vector(20 downto 0);
          Y : in  std_logic_vector(20 downto 0);
          Cin : in  std_logic;
          R : out  std_logic_vector(20 downto 0)   );
end entity;

architecture arch of IntAdder_21_Freq500_uid99 is
signal Rtmp :  std_logic_vector(20 downto 0);
   -- timing of Rtmp: (c17, 0.969231ns)
signal X_d1 :  std_logic_vector(20 downto 0);
   -- timing of X: (c16, 1.569231ns)
signal Y_d1 :  std_logic_vector(20 downto 0);
   -- timing of Y: (c16, 1.569231ns)
signal Cin_d1, Cin_d2, Cin_d3, Cin_d4, Cin_d5, Cin_d6, Cin_d7, Cin_d8, Cin_d9, Cin_d10, Cin_d11, Cin_d12, Cin_d13, Cin_d14, Cin_d15, Cin_d16, Cin_d17 :  std_logic;
   -- timing of Cin: (c0, 0.000000ns)
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            X_d1 <=  X;
            Y_d1 <=  Y;
            Cin_d1 <=  Cin;
            Cin_d2 <=  Cin_d1;
            Cin_d3 <=  Cin_d2;
            Cin_d4 <=  Cin_d3;
            Cin_d5 <=  Cin_d4;
            Cin_d6 <=  Cin_d5;
            Cin_d7 <=  Cin_d6;
            Cin_d8 <=  Cin_d7;
            Cin_d9 <=  Cin_d8;
            Cin_d10 <=  Cin_d9;
            Cin_d11 <=  Cin_d10;
            Cin_d12 <=  Cin_d11;
            Cin_d13 <=  Cin_d12;
            Cin_d14 <=  Cin_d13;
            Cin_d15 <=  Cin_d14;
            Cin_d16 <=  Cin_d15;
            Cin_d17 <=  Cin_d16;
         end if;
      end process;
   Rtmp <= X_d1 + Y_d1 + Cin_d17;
   R <= Rtmp;
end architecture;

--------------------------------------------------------------------------------
--                          FixRealKCM_Freq500_uid89
-- VHDL generated for DummyFPGA @ 500MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin (2007-2016)
--------------------------------------------------------------------------------
-- Pipeline depth: 1 cycles
-- Clock period (ns): 2
-- Target frequency (MHz): 500
-- Input signals: X
-- Output signals: R
--  approx. input signal timings: X: (c16, 1.019231ns)
--  approx. output signal timings: R: (c17, 0.969231ns)

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity FixRealKCM_Freq500_uid89 is
    port (clk : in std_logic;
          X : in  std_logic_vector(7 downto 0);
          R : out  std_logic_vector(20 downto 0)   );
end entity;

architecture arch of FixRealKCM_Freq500_uid89 is
   component FixRealKCM_Freq500_uid89_T0_Freq500_uid92 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(20 downto 0)   );
   end component;

   component FixRealKCM_Freq500_uid89_T1_Freq500_uid95 is
      port ( X : in  std_logic_vector(2 downto 0);
             Y : out  std_logic_vector(15 downto 0)   );
   end component;

   component IntAdder_21_Freq500_uid99 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(20 downto 0);
             Y : in  std_logic_vector(20 downto 0);
             Cin : in  std_logic;
             R : out  std_logic_vector(20 downto 0)   );
   end component;

signal FixRealKCM_Freq500_uid89_A0 :  std_logic_vector(4 downto 0);
   -- timing of FixRealKCM_Freq500_uid89_A0: (c16, 1.019231ns)
signal FixRealKCM_Freq500_uid89_T0 :  std_logic_vector(20 downto 0);
   -- timing of FixRealKCM_Freq500_uid89_T0: (c16, 1.569231ns)
signal FixRealKCM_Freq500_uid89_T0_copy93 :  std_logic_vector(20 downto 0);
   -- timing of FixRealKCM_Freq500_uid89_T0_copy93: (c16, 1.019231ns)
signal bh90_w0_0 :  std_logic;
   -- timing of bh90_w0_0: (c16, 1.569231ns)
signal bh90_w1_0 :  std_logic;
   -- timing of bh90_w1_0: (c16, 1.569231ns)
signal bh90_w2_0 :  std_logic;
   -- timing of bh90_w2_0: (c16, 1.569231ns)
signal bh90_w3_0 :  std_logic;
   -- timing of bh90_w3_0: (c16, 1.569231ns)
signal bh90_w4_0 :  std_logic;
   -- timing of bh90_w4_0: (c16, 1.569231ns)
signal bh90_w5_0 :  std_logic;
   -- timing of bh90_w5_0: (c16, 1.569231ns)
signal bh90_w6_0 :  std_logic;
   -- timing of bh90_w6_0: (c16, 1.569231ns)
signal bh90_w7_0 :  std_logic;
   -- timing of bh90_w7_0: (c16, 1.569231ns)
signal bh90_w8_0 :  std_logic;
   -- timing of bh90_w8_0: (c16, 1.569231ns)
signal bh90_w9_0 :  std_logic;
   -- timing of bh90_w9_0: (c16, 1.569231ns)
signal bh90_w10_0 :  std_logic;
   -- timing of bh90_w10_0: (c16, 1.569231ns)
signal bh90_w11_0 :  std_logic;
   -- timing of bh90_w11_0: (c16, 1.569231ns)
signal bh90_w12_0 :  std_logic;
   -- timing of bh90_w12_0: (c16, 1.569231ns)
signal bh90_w13_0 :  std_logic;
   -- timing of bh90_w13_0: (c16, 1.569231ns)
signal bh90_w14_0 :  std_logic;
   -- timing of bh90_w14_0: (c16, 1.569231ns)
signal bh90_w15_0 :  std_logic;
   -- timing of bh90_w15_0: (c16, 1.569231ns)
signal bh90_w16_0 :  std_logic;
   -- timing of bh90_w16_0: (c16, 1.569231ns)
signal bh90_w17_0 :  std_logic;
   -- timing of bh90_w17_0: (c16, 1.569231ns)
signal bh90_w18_0 :  std_logic;
   -- timing of bh90_w18_0: (c16, 1.569231ns)
signal bh90_w19_0 :  std_logic;
   -- timing of bh90_w19_0: (c16, 1.569231ns)
signal bh90_w20_0 :  std_logic;
   -- timing of bh90_w20_0: (c16, 1.569231ns)
signal FixRealKCM_Freq500_uid89_A1 :  std_logic_vector(2 downto 0);
   -- timing of FixRealKCM_Freq500_uid89_A1: (c16, 1.019231ns)
signal FixRealKCM_Freq500_uid89_T1 :  std_logic_vector(15 downto 0);
   -- timing of FixRealKCM_Freq500_uid89_T1: (c16, 1.569231ns)
signal FixRealKCM_Freq500_uid89_T1_copy96 :  std_logic_vector(15 downto 0);
   -- timing of FixRealKCM_Freq500_uid89_T1_copy96: (c16, 1.019231ns)
signal bh90_w0_1 :  std_logic;
   -- timing of bh90_w0_1: (c16, 1.569231ns)
signal bh90_w1_1 :  std_logic;
   -- timing of bh90_w1_1: (c16, 1.569231ns)
signal bh90_w2_1 :  std_logic;
   -- timing of bh90_w2_1: (c16, 1.569231ns)
signal bh90_w3_1 :  std_logic;
   -- timing of bh90_w3_1: (c16, 1.569231ns)
signal bh90_w4_1 :  std_logic;
   -- timing of bh90_w4_1: (c16, 1.569231ns)
signal bh90_w5_1 :  std_logic;
   -- timing of bh90_w5_1: (c16, 1.569231ns)
signal bh90_w6_1 :  std_logic;
   -- timing of bh90_w6_1: (c16, 1.569231ns)
signal bh90_w7_1 :  std_logic;
   -- timing of bh90_w7_1: (c16, 1.569231ns)
signal bh90_w8_1 :  std_logic;
   -- timing of bh90_w8_1: (c16, 1.569231ns)
signal bh90_w9_1 :  std_logic;
   -- timing of bh90_w9_1: (c16, 1.569231ns)
signal bh90_w10_1 :  std_logic;
   -- timing of bh90_w10_1: (c16, 1.569231ns)
signal bh90_w11_1 :  std_logic;
   -- timing of bh90_w11_1: (c16, 1.569231ns)
signal bh90_w12_1 :  std_logic;
   -- timing of bh90_w12_1: (c16, 1.569231ns)
signal bh90_w13_1 :  std_logic;
   -- timing of bh90_w13_1: (c16, 1.569231ns)
signal bh90_w14_1 :  std_logic;
   -- timing of bh90_w14_1: (c16, 1.569231ns)
signal bh90_w15_1 :  std_logic;
   -- timing of bh90_w15_1: (c16, 1.569231ns)
signal bitheapFinalAdd_bh90_In0 :  std_logic_vector(20 downto 0);
   -- timing of bitheapFinalAdd_bh90_In0: (c16, 1.569231ns)
signal bitheapFinalAdd_bh90_In1 :  std_logic_vector(20 downto 0);
   -- timing of bitheapFinalAdd_bh90_In1: (c16, 1.569231ns)
signal bitheapFinalAdd_bh90_Cin :  std_logic;
   -- timing of bitheapFinalAdd_bh90_Cin: (c0, 0.000000ns)
signal bitheapFinalAdd_bh90_Out :  std_logic_vector(20 downto 0);
   -- timing of bitheapFinalAdd_bh90_Out: (c17, 0.969231ns)
signal bitheapResult_bh90 :  std_logic_vector(20 downto 0);
   -- timing of bitheapResult_bh90: (c17, 0.969231ns)
signal OutRes :  std_logic_vector(20 downto 0);
   -- timing of OutRes: (c17, 0.969231ns)
begin
-- This operator multiplies by log(2)
   FixRealKCM_Freq500_uid89_A0 <= X(7 downto 3);-- input address  m=7  l=3
   FixRealKCM_Freq500_uid89_Table0: FixRealKCM_Freq500_uid89_T0_Freq500_uid92
      port map ( X => FixRealKCM_Freq500_uid89_A0,
                 Y => FixRealKCM_Freq500_uid89_T0_copy93);
   FixRealKCM_Freq500_uid89_T0 <= FixRealKCM_Freq500_uid89_T0_copy93; -- output copy to hold a pipeline register if needed
   bh90_w0_0 <= FixRealKCM_Freq500_uid89_T0(0);
   bh90_w1_0 <= FixRealKCM_Freq500_uid89_T0(1);
   bh90_w2_0 <= FixRealKCM_Freq500_uid89_T0(2);
   bh90_w3_0 <= FixRealKCM_Freq500_uid89_T0(3);
   bh90_w4_0 <= FixRealKCM_Freq500_uid89_T0(4);
   bh90_w5_0 <= FixRealKCM_Freq500_uid89_T0(5);
   bh90_w6_0 <= FixRealKCM_Freq500_uid89_T0(6);
   bh90_w7_0 <= FixRealKCM_Freq500_uid89_T0(7);
   bh90_w8_0 <= FixRealKCM_Freq500_uid89_T0(8);
   bh90_w9_0 <= FixRealKCM_Freq500_uid89_T0(9);
   bh90_w10_0 <= FixRealKCM_Freq500_uid89_T0(10);
   bh90_w11_0 <= FixRealKCM_Freq500_uid89_T0(11);
   bh90_w12_0 <= FixRealKCM_Freq500_uid89_T0(12);
   bh90_w13_0 <= FixRealKCM_Freq500_uid89_T0(13);
   bh90_w14_0 <= FixRealKCM_Freq500_uid89_T0(14);
   bh90_w15_0 <= FixRealKCM_Freq500_uid89_T0(15);
   bh90_w16_0 <= FixRealKCM_Freq500_uid89_T0(16);
   bh90_w17_0 <= FixRealKCM_Freq500_uid89_T0(17);
   bh90_w18_0 <= FixRealKCM_Freq500_uid89_T0(18);
   bh90_w19_0 <= FixRealKCM_Freq500_uid89_T0(19);
   bh90_w20_0 <= FixRealKCM_Freq500_uid89_T0(20);
   FixRealKCM_Freq500_uid89_A1 <= X(2 downto 0);-- input address  m=2  l=0
   FixRealKCM_Freq500_uid89_Table1: FixRealKCM_Freq500_uid89_T1_Freq500_uid95
      port map ( X => FixRealKCM_Freq500_uid89_A1,
                 Y => FixRealKCM_Freq500_uid89_T1_copy96);
   FixRealKCM_Freq500_uid89_T1 <= FixRealKCM_Freq500_uid89_T1_copy96; -- output copy to hold a pipeline register if needed
   bh90_w0_1 <= FixRealKCM_Freq500_uid89_T1(0);
   bh90_w1_1 <= FixRealKCM_Freq500_uid89_T1(1);
   bh90_w2_1 <= FixRealKCM_Freq500_uid89_T1(2);
   bh90_w3_1 <= FixRealKCM_Freq500_uid89_T1(3);
   bh90_w4_1 <= FixRealKCM_Freq500_uid89_T1(4);
   bh90_w5_1 <= FixRealKCM_Freq500_uid89_T1(5);
   bh90_w6_1 <= FixRealKCM_Freq500_uid89_T1(6);
   bh90_w7_1 <= FixRealKCM_Freq500_uid89_T1(7);
   bh90_w8_1 <= FixRealKCM_Freq500_uid89_T1(8);
   bh90_w9_1 <= FixRealKCM_Freq500_uid89_T1(9);
   bh90_w10_1 <= FixRealKCM_Freq500_uid89_T1(10);
   bh90_w11_1 <= FixRealKCM_Freq500_uid89_T1(11);
   bh90_w12_1 <= FixRealKCM_Freq500_uid89_T1(12);
   bh90_w13_1 <= FixRealKCM_Freq500_uid89_T1(13);
   bh90_w14_1 <= FixRealKCM_Freq500_uid89_T1(14);
   bh90_w15_1 <= FixRealKCM_Freq500_uid89_T1(15);

   -- Adding the constant bits 
      -- All the constant bits are zero, nothing to add


   bitheapFinalAdd_bh90_In0 <= "" & bh90_w20_0 & bh90_w19_0 & bh90_w18_0 & bh90_w17_0 & bh90_w16_0 & bh90_w15_0 & bh90_w14_0 & bh90_w13_0 & bh90_w12_0 & bh90_w11_0 & bh90_w10_0 & bh90_w9_0 & bh90_w8_0 & bh90_w7_0 & bh90_w6_0 & bh90_w5_0 & bh90_w4_0 & bh90_w3_0 & bh90_w2_0 & bh90_w1_0 & bh90_w0_0;
   bitheapFinalAdd_bh90_In1 <= "0" & "0" & "0" & "0" & "0" & bh90_w15_1 & bh90_w14_1 & bh90_w13_1 & bh90_w12_1 & bh90_w11_1 & bh90_w10_1 & bh90_w9_1 & bh90_w8_1 & bh90_w7_1 & bh90_w6_1 & bh90_w5_1 & bh90_w4_1 & bh90_w3_1 & bh90_w2_1 & bh90_w1_1 & bh90_w0_1;
   bitheapFinalAdd_bh90_Cin <= '0';

   bitheapFinalAdd_bh90: IntAdder_21_Freq500_uid99
      port map ( clk  => clk,
                 Cin => bitheapFinalAdd_bh90_Cin,
                 X => bitheapFinalAdd_bh90_In0,
                 Y => bitheapFinalAdd_bh90_In1,
                 R => bitheapFinalAdd_bh90_Out);
   bitheapResult_bh90 <= bitheapFinalAdd_bh90_Out(20 downto 0);
   OutRes <= bitheapResult_bh90(20 downto 0);
   R <= OutRes(20 downto 0);
end architecture;

--------------------------------------------------------------------------------
--                         IntAdder_13_Freq500_uid102
-- VHDL generated for DummyFPGA @ 500MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin (2008-2016)
--------------------------------------------------------------------------------
-- Pipeline depth: 18 cycles
-- Clock period (ns): 2
-- Target frequency (MHz): 500
-- Input signals: X Y Cin
-- Output signals: R
--  approx. input signal timings: X: (c15, 1.709231ns)Y: (c17, 0.969231ns)Cin: (c0, 0.000000ns)
--  approx. output signal timings: R: (c18, 0.289231ns)

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntAdder_13_Freq500_uid102 is
    port (clk : in std_logic;
          X : in  std_logic_vector(12 downto 0);
          Y : in  std_logic_vector(12 downto 0);
          Cin : in  std_logic;
          R : out  std_logic_vector(12 downto 0)   );
end entity;

architecture arch of IntAdder_13_Freq500_uid102 is
signal Rtmp :  std_logic_vector(12 downto 0);
   -- timing of Rtmp: (c18, 0.289231ns)
signal X_d1, X_d2, X_d3 :  std_logic_vector(12 downto 0);
   -- timing of X: (c15, 1.709231ns)
signal Y_d1 :  std_logic_vector(12 downto 0);
   -- timing of Y: (c17, 0.969231ns)
signal Cin_d1, Cin_d2, Cin_d3, Cin_d4, Cin_d5, Cin_d6, Cin_d7, Cin_d8, Cin_d9, Cin_d10, Cin_d11, Cin_d12, Cin_d13, Cin_d14, Cin_d15, Cin_d16, Cin_d17, Cin_d18 :  std_logic;
   -- timing of Cin: (c0, 0.000000ns)
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            X_d1 <=  X;
            X_d2 <=  X_d1;
            X_d3 <=  X_d2;
            Y_d1 <=  Y;
            Cin_d1 <=  Cin;
            Cin_d2 <=  Cin_d1;
            Cin_d3 <=  Cin_d2;
            Cin_d4 <=  Cin_d3;
            Cin_d5 <=  Cin_d4;
            Cin_d6 <=  Cin_d5;
            Cin_d7 <=  Cin_d6;
            Cin_d8 <=  Cin_d7;
            Cin_d9 <=  Cin_d8;
            Cin_d10 <=  Cin_d9;
            Cin_d11 <=  Cin_d10;
            Cin_d12 <=  Cin_d11;
            Cin_d13 <=  Cin_d12;
            Cin_d14 <=  Cin_d13;
            Cin_d15 <=  Cin_d14;
            Cin_d16 <=  Cin_d15;
            Cin_d17 <=  Cin_d16;
            Cin_d18 <=  Cin_d17;
         end if;
      end process;
   Rtmp <= X_d3 + Y_d1 + Cin_d18;
   R <= Rtmp;
end architecture;

--------------------------------------------------------------------------------
--                         IntAdder_4_Freq500_uid112
-- VHDL generated for DummyFPGA @ 500MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin (2008-2016)
--------------------------------------------------------------------------------
-- Pipeline depth: 19 cycles
-- Clock period (ns): 2
-- Target frequency (MHz): 500
-- Input signals: X Y Cin
-- Output signals: R
--  approx. input signal timings: X: (c18, 0.839231ns)Y: (c0, 0.000000ns)Cin: (c0, 0.000000ns)
--  approx. output signal timings: R: (c19, 0.069231ns)

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntAdder_4_Freq500_uid112 is
    port (clk : in std_logic;
          X : in  std_logic_vector(3 downto 0);
          Y : in  std_logic_vector(3 downto 0);
          Cin : in  std_logic;
          R : out  std_logic_vector(3 downto 0)   );
end entity;

architecture arch of IntAdder_4_Freq500_uid112 is
signal Rtmp :  std_logic_vector(3 downto 0);
   -- timing of Rtmp: (c19, 0.069231ns)
signal X_d1 :  std_logic_vector(3 downto 0);
   -- timing of X: (c18, 0.839231ns)
signal Y_d1, Y_d2, Y_d3, Y_d4, Y_d5, Y_d6, Y_d7, Y_d8, Y_d9, Y_d10, Y_d11, Y_d12, Y_d13, Y_d14, Y_d15, Y_d16, Y_d17, Y_d18, Y_d19 :  std_logic_vector(3 downto 0);
   -- timing of Y: (c0, 0.000000ns)
signal Cin_d1, Cin_d2, Cin_d3, Cin_d4, Cin_d5, Cin_d6, Cin_d7, Cin_d8, Cin_d9, Cin_d10, Cin_d11, Cin_d12, Cin_d13, Cin_d14, Cin_d15, Cin_d16, Cin_d17, Cin_d18, Cin_d19 :  std_logic;
   -- timing of Cin: (c0, 0.000000ns)
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            X_d1 <=  X;
            Y_d1 <=  Y;
            Y_d2 <=  Y_d1;
            Y_d3 <=  Y_d2;
            Y_d4 <=  Y_d3;
            Y_d5 <=  Y_d4;
            Y_d6 <=  Y_d5;
            Y_d7 <=  Y_d6;
            Y_d8 <=  Y_d7;
            Y_d9 <=  Y_d8;
            Y_d10 <=  Y_d9;
            Y_d11 <=  Y_d10;
            Y_d12 <=  Y_d11;
            Y_d13 <=  Y_d12;
            Y_d14 <=  Y_d13;
            Y_d15 <=  Y_d14;
            Y_d16 <=  Y_d15;
            Y_d17 <=  Y_d16;
            Y_d18 <=  Y_d17;
            Y_d19 <=  Y_d18;
            Cin_d1 <=  Cin;
            Cin_d2 <=  Cin_d1;
            Cin_d3 <=  Cin_d2;
            Cin_d4 <=  Cin_d3;
            Cin_d5 <=  Cin_d4;
            Cin_d6 <=  Cin_d5;
            Cin_d7 <=  Cin_d6;
            Cin_d8 <=  Cin_d7;
            Cin_d9 <=  Cin_d8;
            Cin_d10 <=  Cin_d9;
            Cin_d11 <=  Cin_d10;
            Cin_d12 <=  Cin_d11;
            Cin_d13 <=  Cin_d12;
            Cin_d14 <=  Cin_d13;
            Cin_d15 <=  Cin_d14;
            Cin_d16 <=  Cin_d15;
            Cin_d17 <=  Cin_d16;
            Cin_d18 <=  Cin_d17;
            Cin_d19 <=  Cin_d18;
         end if;
      end process;
   Rtmp <= X_d1 + Y_d19 + Cin_d19;
   R <= Rtmp;
end architecture;

--------------------------------------------------------------------------------
--                     IntMultiplier_3x4_5_Freq500_uid114
-- VHDL generated for DummyFPGA @ 500MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Martin Kumm, Florent de Dinechin, Andreas Böttcher, Kinga Illyes, Bogdan Popa, Bogdan Pasca, 2012-
--------------------------------------------------------------------------------
-- Pipeline depth: 1 cycles
-- Clock period (ns): 2
-- Target frequency (MHz): 500
-- Input signals: X Y
-- Output signals: R
--  approx. input signal timings: X: (c19, 0.069231ns)Y: (c18, 0.839231ns)
--  approx. output signal timings: R: (c19, 0.069231ns)

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity IntMultiplier_3x4_5_Freq500_uid114 is
    port (clk : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(3 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplier_3x4_5_Freq500_uid114 is
signal XX_m115 :  std_logic_vector(2 downto 0);
   -- timing of XX_m115: (c19, 0.069231ns)
signal YY_m115 :  std_logic_vector(3 downto 0);
   -- timing of YY_m115: (c18, 0.839231ns)
signal XX :  unsigned(-1+3 downto 0);
   -- timing of XX: (c19, 0.069231ns)
signal YY, YY_d1 :  unsigned(-1+4 downto 0);
   -- timing of YY: (c18, 0.839231ns)
signal RR :  unsigned(-1+7 downto 0);
   -- timing of RR: (c19, 0.069231ns)
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            YY_d1 <=  YY;
         end if;
      end process;
   XX_m115 <= X ;
   YY_m115 <= Y ;
   XX <= unsigned(X);
   YY <= unsigned(Y);
   RR <= XX*YY_d1;
   R <= std_logic_vector(RR(6 downto 2));
end architecture;

--------------------------------------------------------------------------------
--                         IntAdder_14_Freq500_uid118
-- VHDL generated for DummyFPGA @ 500MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin (2008-2016)
--------------------------------------------------------------------------------
-- Pipeline depth: 19 cycles
-- Clock period (ns): 2
-- Target frequency (MHz): 500
-- Input signals: X Y Cin
-- Output signals: R
--  approx. input signal timings: X: (c18, 0.839231ns)Y: (c19, 0.069231ns)Cin: (c0, 0.000000ns)
--  approx. output signal timings: R: (c19, 1.199231ns)

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntAdder_14_Freq500_uid118 is
    port (clk : in std_logic;
          X : in  std_logic_vector(13 downto 0);
          Y : in  std_logic_vector(13 downto 0);
          Cin : in  std_logic;
          R : out  std_logic_vector(13 downto 0)   );
end entity;

architecture arch of IntAdder_14_Freq500_uid118 is
signal Rtmp :  std_logic_vector(13 downto 0);
   -- timing of Rtmp: (c19, 1.199231ns)
signal X_d1 :  std_logic_vector(13 downto 0);
   -- timing of X: (c18, 0.839231ns)
signal Cin_d1, Cin_d2, Cin_d3, Cin_d4, Cin_d5, Cin_d6, Cin_d7, Cin_d8, Cin_d9, Cin_d10, Cin_d11, Cin_d12, Cin_d13, Cin_d14, Cin_d15, Cin_d16, Cin_d17, Cin_d18, Cin_d19 :  std_logic;
   -- timing of Cin: (c0, 0.000000ns)
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            X_d1 <=  X;
            Cin_d1 <=  Cin;
            Cin_d2 <=  Cin_d1;
            Cin_d3 <=  Cin_d2;
            Cin_d4 <=  Cin_d3;
            Cin_d5 <=  Cin_d4;
            Cin_d6 <=  Cin_d5;
            Cin_d7 <=  Cin_d6;
            Cin_d8 <=  Cin_d7;
            Cin_d9 <=  Cin_d8;
            Cin_d10 <=  Cin_d9;
            Cin_d11 <=  Cin_d10;
            Cin_d12 <=  Cin_d11;
            Cin_d13 <=  Cin_d12;
            Cin_d14 <=  Cin_d13;
            Cin_d15 <=  Cin_d14;
            Cin_d16 <=  Cin_d15;
            Cin_d17 <=  Cin_d16;
            Cin_d18 <=  Cin_d17;
            Cin_d19 <=  Cin_d18;
         end if;
      end process;
   Rtmp <= X_d1 + Y + Cin_d19;
   R <= Rtmp;
end architecture;

--------------------------------------------------------------------------------
--                           Exp_8_10_Freq500_uid75
-- VHDL generated for DummyFPGA @ 500MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: F. de Dinechin, Bogdan Pasca, Orégane Desrentes (2008-2025)
--------------------------------------------------------------------------------
-- Pipeline depth: 6 cycles
-- Clock period (ns): 2
-- Target frequency (MHz): 500
-- Input signals: ufixX_i XSign
-- Output signals: expY K
--  approx. input signal timings: ufixX_i: (c15, 1.159231ns)XSign: (c13, 1.615385ns)
--  approx. output signal timings: expY: (c19, 1.199231ns)K: (c17, 0.299231ns)

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity Exp_8_10_Freq500_uid75 is
    port (clk : in std_logic;
          ufixX_i : in  std_logic_vector(19 downto 0);
          XSign : in  std_logic;
          expY : out  std_logic_vector(13 downto 0);
          K : out  std_logic_vector(8 downto 0)   );
end entity;

architecture arch of Exp_8_10_Freq500_uid75 is
   component FixRealKCM_Freq500_uid77 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(9 downto 0);
             R : out  std_logic_vector(7 downto 0)   );
   end component;

   component FixRealKCM_Freq500_uid89 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(7 downto 0);
             R : out  std_logic_vector(20 downto 0)   );
   end component;

   component IntAdder_13_Freq500_uid102 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(12 downto 0);
             Y : in  std_logic_vector(12 downto 0);
             Cin : in  std_logic;
             R : out  std_logic_vector(12 downto 0)   );
   end component;

   component FixFunctionByTable_Freq500_uid104 is
      port ( X : in  std_logic_vector(9 downto 0);
             Y : out  std_logic_vector(13 downto 0)   );
   end component;

   component FixFunctionByTable_Freq500_uid107 is
      port ( X : in  std_logic_vector(2 downto 0);
             Y : out  std_logic_vector(2 downto 0)   );
   end component;

   component IntAdder_4_Freq500_uid112 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(3 downto 0);
             Y : in  std_logic_vector(3 downto 0);
             Cin : in  std_logic;
             R : out  std_logic_vector(3 downto 0)   );
   end component;

   component IntMultiplier_3x4_5_Freq500_uid114 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(3 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntAdder_14_Freq500_uid118 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(13 downto 0);
             Y : in  std_logic_vector(13 downto 0);
             Cin : in  std_logic;
             R : out  std_logic_vector(13 downto 0)   );
   end component;

signal ufixX :  unsigned(6+13 downto 0);
   -- timing of ufixX: (c15, 1.159231ns)
signal xMulIn :  unsigned(6+3 downto 0);
   -- timing of xMulIn: (c15, 1.159231ns)
signal absK, absK_d1 :  std_logic_vector(7 downto 0);
   -- timing of absK: (c16, 1.019231ns)
signal minusAbsK :  std_logic_vector(8 downto 0);
   -- timing of minusAbsK: (c17, 0.299231ns)
signal absKLog2 :  std_logic_vector(20 downto 0);
   -- timing of absKLog2: (c17, 0.969231ns)
signal subOp1 :  std_logic_vector(12 downto 0);
   -- timing of subOp1: (c15, 1.709231ns)
signal subOp2 :  std_logic_vector(12 downto 0);
   -- timing of subOp2: (c17, 0.969231ns)
signal Y :  std_logic_vector(12 downto 0);
   -- timing of Y: (c18, 0.289231ns)
signal A :  std_logic_vector(9 downto 0);
   -- timing of A: (c18, 0.289231ns)
signal Z :  std_logic_vector(2 downto 0);
   -- timing of Z: (c18, 0.289231ns)
signal expA :  std_logic_vector(13 downto 0);
   -- timing of expA: (c18, 0.839231ns)
signal expA_copy105 :  std_logic_vector(13 downto 0);
   -- timing of expA_copy105: (c18, 0.289231ns)
signal expZm1_p :  std_logic_vector(2 downto 0);
   -- timing of expZm1_p: (c18, 0.839231ns)
signal expZm1_p_copy108 :  std_logic_vector(2 downto 0);
   -- timing of expZm1_p_copy108: (c18, 0.289231ns)
signal expZm1 :  std_logic_vector(3 downto 0);
   -- timing of expZm1: (c18, 0.839231ns)
signal expA_T :  std_logic_vector(3 downto 0);
   -- timing of expA_T: (c18, 0.839231ns)
signal expArounded0 :  std_logic_vector(3 downto 0);
   -- timing of expArounded0: (c19, 0.069231ns)
signal expArounded :  std_logic_vector(2 downto 0);
   -- timing of expArounded: (c19, 0.069231ns)
signal lowerProduct :  std_logic_vector(4 downto 0);
   -- timing of lowerProduct: (c19, 0.069231ns)
signal extendedLowerProduct :  std_logic_vector(13 downto 0);
   -- timing of extendedLowerProduct: (c19, 0.069231ns)
signal XSign_d1, XSign_d2, XSign_d3, XSign_d4 :  std_logic;
   -- timing of XSign: (c13, 1.615385ns)
constant g: positive := 3;
constant wE: positive := 8;
constant wF: positive := 10;
constant wFIn: positive := 10;
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            absK_d1 <=  absK;
            XSign_d1 <=  XSign;
            XSign_d2 <=  XSign_d1;
            XSign_d3 <=  XSign_d2;
            XSign_d4 <=  XSign_d3;
         end if;
      end process;
ufixX <= unsigned(ufixX_i);
   xMulIn <= ufixX(19 downto 10); -- fix resize from (6, -13) to (6, -3)
   MulInvLog2: FixRealKCM_Freq500_uid77
      port map ( clk  => clk,
                 X => std_logic_vector(xMulIn),
                 R => absK);
   minusAbsK <= (8 downto 0 => '0') - ('0' & absK_d1);
   K <= minusAbsK when  XSign_d4='1'   else ('0' & absK_d1);
   MulLog2: FixRealKCM_Freq500_uid89
      port map ( clk  => clk,
                 X => absK,
                 R => absKLog2);
   subOp1 <= std_logic_vector(ufixX(12 downto 0)) when XSign_d2='0' else not (std_logic_vector(ufixX(12 downto 0)));
   subOp2 <= absKLog2(12 downto 0) when XSign_d4='1' else not (absKLog2(12 downto 0));
   theYAdder: IntAdder_13_Freq500_uid102
      port map ( clk  => clk,
                 Cin => '1',
                 X => subOp1,
                 Y => subOp2,
                 R => Y);
   -- Now compute the exp of this fixed-point value
   A <= Y(12 downto 3);
   Z <= Y(2 downto 0);
   ExpATable: FixFunctionByTable_Freq500_uid104
      port map ( X => A,
                 Y => expA_copy105);
   expA <= expA_copy105; -- output copy to hold a pipeline register if needed
   ExpZm1Table: FixFunctionByTable_Freq500_uid107
      port map ( X => Z,
                 Y => expZm1_p_copy108);
   expZm1_p <= expZm1_p_copy108; -- output copy to hold a pipeline register if needed
expZm1 <= "0" & expZm1_p;
   -- Rounding expA to the same accuracy as expZm1
   --   (truncation would not be accurate enough and require one more guard bit)
   expA_T <= expA(13 downto 10);
   Adder_expArounded0: IntAdder_4_Freq500_uid112
      port map ( clk  => clk,
                 Cin => '1',
                 X => expA_T,
                 Y => "0000",
                 R => expArounded0);
   expArounded <= expArounded0(3 downto 1);
   TheLowerProduct: IntMultiplier_3x4_5_Freq500_uid114
      port map ( clk  => clk,
                 X => expArounded,
                 Y => expZm1,
                 R => lowerProduct);
   extendedLowerProduct <= ((13 downto 5 => '0') & lowerProduct(4 downto 0));
   -- Final addition -- the product MSB bit weight is -k+2 = -8
   TheFinalAdder: IntAdder_14_Freq500_uid118
      port map ( clk  => clk,
                 Cin => '0',
                 X => expA,
                 Y => extendedLowerProduct,
                 R => expY);
end architecture;

--------------------------------------------------------------------------------
--                         IntAdder_20_Freq500_uid121
-- VHDL generated for DummyFPGA @ 500MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin (2008-2016)
--------------------------------------------------------------------------------
-- Pipeline depth: 20 cycles
-- Clock period (ns): 2
-- Target frequency (MHz): 500
-- Input signals: X Y Cin
-- Output signals: R
--  approx. input signal timings: X: (c19, 1.749231ns)Y: (c19, 1.199231ns)Cin: (c0, 0.000000ns)
--  approx. output signal timings: R: (c20, 1.139231ns)

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntAdder_20_Freq500_uid121 is
    port (clk : in std_logic;
          X : in  std_logic_vector(19 downto 0);
          Y : in  std_logic_vector(19 downto 0);
          Cin : in  std_logic;
          R : out  std_logic_vector(19 downto 0)   );
end entity;

architecture arch of IntAdder_20_Freq500_uid121 is
signal Rtmp :  std_logic_vector(19 downto 0);
   -- timing of Rtmp: (c20, 1.139231ns)
signal X_d1 :  std_logic_vector(19 downto 0);
   -- timing of X: (c19, 1.749231ns)
signal Y_d1 :  std_logic_vector(19 downto 0);
   -- timing of Y: (c19, 1.199231ns)
signal Cin_d1, Cin_d2, Cin_d3, Cin_d4, Cin_d5, Cin_d6, Cin_d7, Cin_d8, Cin_d9, Cin_d10, Cin_d11, Cin_d12, Cin_d13, Cin_d14, Cin_d15, Cin_d16, Cin_d17, Cin_d18, Cin_d19, Cin_d20 :  std_logic;
   -- timing of Cin: (c0, 0.000000ns)
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            X_d1 <=  X;
            Y_d1 <=  Y;
            Cin_d1 <=  Cin;
            Cin_d2 <=  Cin_d1;
            Cin_d3 <=  Cin_d2;
            Cin_d4 <=  Cin_d3;
            Cin_d5 <=  Cin_d4;
            Cin_d6 <=  Cin_d5;
            Cin_d7 <=  Cin_d6;
            Cin_d8 <=  Cin_d7;
            Cin_d9 <=  Cin_d8;
            Cin_d10 <=  Cin_d9;
            Cin_d11 <=  Cin_d10;
            Cin_d12 <=  Cin_d11;
            Cin_d13 <=  Cin_d12;
            Cin_d14 <=  Cin_d13;
            Cin_d15 <=  Cin_d14;
            Cin_d16 <=  Cin_d15;
            Cin_d17 <=  Cin_d16;
            Cin_d18 <=  Cin_d17;
            Cin_d19 <=  Cin_d18;
            Cin_d20 <=  Cin_d19;
         end if;
      end process;
   Rtmp <= X_d1 + Y_d1 + Cin_d20;
   R <= Rtmp;
end architecture;

--------------------------------------------------------------------------------
--                          FPExp_8_10_Freq500_uid71
-- VHDL generated for DummyFPGA @ 500MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: F. de Dinechin, Bogdan Pasca, Orégane Desrentes (2008-2025)
--------------------------------------------------------------------------------
-- Pipeline depth: 7 cycles
-- Clock period (ns): 2
-- Target frequency (MHz): 500
-- Input signals: X
-- Output signals: R
--  approx. input signal timings: X: (c13, 1.615385ns)
--  approx. output signal timings: R: (c20, 1.689231ns)

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity FPExp_8_10_Freq500_uid71 is
    port (clk : in std_logic;
          X : in  std_logic_vector(8+21+2 downto 0);
          R : out  std_logic_vector(8+10+2 downto 0)   );
end entity;

architecture arch of FPExp_8_10_Freq500_uid71 is
   component LeftShifter22_by_max_19_Freq500_uid73 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(21 downto 0);
             S : in  std_logic_vector(4 downto 0);
             R : out  std_logic_vector(40 downto 0)   );
   end component;

   component Exp_8_10_Freq500_uid75 is
      port ( clk : in std_logic;
             ufixX_i : in  std_logic_vector(19 downto 0);
             XSign : in  std_logic;
             expY : out  std_logic_vector(13 downto 0);
             K : out  std_logic_vector(8 downto 0)   );
   end component;

   component IntAdder_20_Freq500_uid121 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(19 downto 0);
             Y : in  std_logic_vector(19 downto 0);
             Cin : in  std_logic;
             R : out  std_logic_vector(19 downto 0)   );
   end component;

signal Xexn, Xexn_d1, Xexn_d2, Xexn_d3, Xexn_d4, Xexn_d5, Xexn_d6, Xexn_d7 :  std_logic_vector(1 downto 0);
   -- timing of Xexn: (c13, 1.615385ns)
signal XSign, XSign_d1, XSign_d2, XSign_d3, XSign_d4, XSign_d5, XSign_d6, XSign_d7 :  std_logic;
   -- timing of XSign: (c13, 1.615385ns)
signal XexpField, XexpField_d1 :  std_logic_vector(7 downto 0);
   -- timing of XexpField: (c13, 1.615385ns)
signal Xfrac :  unsigned(-1+21 downto 0);
   -- timing of Xfrac: (c13, 1.615385ns)
signal e0, e0_d1, e0_d2, e0_d3, e0_d4, e0_d5, e0_d6, e0_d7, e0_d8, e0_d9, e0_d10, e0_d11, e0_d12, e0_d13, e0_d14 :  std_logic_vector(9 downto 0);
   -- timing of e0: (c0, 0.000000ns)
signal shiftVal, shiftVal_d1 :  std_logic_vector(9 downto 0);
   -- timing of shiftVal: (c14, 0.905385ns)
signal resultWillBeOne, resultWillBeOne_d1 :  std_logic;
   -- timing of resultWillBeOne: (c14, 0.905385ns)
signal mXu :  unsigned(0+21 downto 0);
   -- timing of mXu: (c13, 1.615385ns)
signal maxShift, maxShift_d1, maxShift_d2, maxShift_d3, maxShift_d4, maxShift_d5, maxShift_d6, maxShift_d7, maxShift_d8, maxShift_d9, maxShift_d10, maxShift_d11, maxShift_d12, maxShift_d13, maxShift_d14, maxShift_d15 :  std_logic_vector(8 downto 0);
   -- timing of maxShift: (c0, 0.000000ns)
signal overflow0 :  std_logic;
   -- timing of overflow0: (c15, 0.185385ns)
signal shiftValIn :  std_logic_vector(4 downto 0);
   -- timing of shiftValIn: (c14, 0.905385ns)
signal fixX0 :  std_logic_vector(40 downto 0);
   -- timing of fixX0: (c15, 1.159231ns)
signal ufixX :  unsigned(6+13 downto 0);
   -- timing of ufixX: (c15, 1.159231ns)
signal expY :  std_logic_vector(13 downto 0);
   -- timing of expY: (c19, 1.199231ns)
signal K, K_d1, K_d2 :  std_logic_vector(8 downto 0);
   -- timing of K: (c17, 0.299231ns)
signal needNoNorm :  std_logic;
   -- timing of needNoNorm: (c19, 1.199231ns)
signal preRoundBiasSig :  std_logic_vector(19 downto 0);
   -- timing of preRoundBiasSig: (c19, 1.749231ns)
signal roundBit :  std_logic;
   -- timing of roundBit: (c19, 1.199231ns)
signal roundNormAddend :  std_logic_vector(19 downto 0);
   -- timing of roundNormAddend: (c19, 1.199231ns)
signal roundedExpSigRes :  std_logic_vector(19 downto 0);
   -- timing of roundedExpSigRes: (c20, 1.139231ns)
signal roundedExpSig :  std_logic_vector(19 downto 0);
   -- timing of roundedExpSig: (c20, 1.689231ns)
signal ofl1, ofl1_d1, ofl1_d2, ofl1_d3, ofl1_d4, ofl1_d5 :  std_logic;
   -- timing of ofl1: (c15, 0.735385ns)
signal ofl2 :  std_logic;
   -- timing of ofl2: (c20, 1.689231ns)
signal ofl3, ofl3_d1, ofl3_d2, ofl3_d3, ofl3_d4, ofl3_d5, ofl3_d6, ofl3_d7 :  std_logic;
   -- timing of ofl3: (c13, 1.615385ns)
signal ofl :  std_logic;
   -- timing of ofl: (c20, 1.689231ns)
signal ufl1 :  std_logic;
   -- timing of ufl1: (c20, 1.689231ns)
signal ufl2, ufl2_d1, ufl2_d2, ufl2_d3, ufl2_d4, ufl2_d5, ufl2_d6, ufl2_d7 :  std_logic;
   -- timing of ufl2: (c13, 1.615385ns)
signal ufl3, ufl3_d1, ufl3_d2, ufl3_d3, ufl3_d4, ufl3_d5 :  std_logic;
   -- timing of ufl3: (c15, 0.185385ns)
signal ufl :  std_logic;
   -- timing of ufl: (c20, 1.689231ns)
signal Rexn :  std_logic_vector(1 downto 0);
   -- timing of Rexn: (c20, 1.689231ns)
constant g: positive := 3;
constant wE: positive := 8;
constant wF: positive := 10;
constant wFIn: positive := 21;
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            Xexn_d1 <=  Xexn;
            Xexn_d2 <=  Xexn_d1;
            Xexn_d3 <=  Xexn_d2;
            Xexn_d4 <=  Xexn_d3;
            Xexn_d5 <=  Xexn_d4;
            Xexn_d6 <=  Xexn_d5;
            Xexn_d7 <=  Xexn_d6;
            XSign_d1 <=  XSign;
            XSign_d2 <=  XSign_d1;
            XSign_d3 <=  XSign_d2;
            XSign_d4 <=  XSign_d3;
            XSign_d5 <=  XSign_d4;
            XSign_d6 <=  XSign_d5;
            XSign_d7 <=  XSign_d6;
            XexpField_d1 <=  XexpField;
            e0_d1 <=  e0;
            e0_d2 <=  e0_d1;
            e0_d3 <=  e0_d2;
            e0_d4 <=  e0_d3;
            e0_d5 <=  e0_d4;
            e0_d6 <=  e0_d5;
            e0_d7 <=  e0_d6;
            e0_d8 <=  e0_d7;
            e0_d9 <=  e0_d8;
            e0_d10 <=  e0_d9;
            e0_d11 <=  e0_d10;
            e0_d12 <=  e0_d11;
            e0_d13 <=  e0_d12;
            e0_d14 <=  e0_d13;
            shiftVal_d1 <=  shiftVal;
            resultWillBeOne_d1 <=  resultWillBeOne;
            maxShift_d1 <=  maxShift;
            maxShift_d2 <=  maxShift_d1;
            maxShift_d3 <=  maxShift_d2;
            maxShift_d4 <=  maxShift_d3;
            maxShift_d5 <=  maxShift_d4;
            maxShift_d6 <=  maxShift_d5;
            maxShift_d7 <=  maxShift_d6;
            maxShift_d8 <=  maxShift_d7;
            maxShift_d9 <=  maxShift_d8;
            maxShift_d10 <=  maxShift_d9;
            maxShift_d11 <=  maxShift_d10;
            maxShift_d12 <=  maxShift_d11;
            maxShift_d13 <=  maxShift_d12;
            maxShift_d14 <=  maxShift_d13;
            maxShift_d15 <=  maxShift_d14;
            K_d1 <=  K;
            K_d2 <=  K_d1;
            ofl1_d1 <=  ofl1;
            ofl1_d2 <=  ofl1_d1;
            ofl1_d3 <=  ofl1_d2;
            ofl1_d4 <=  ofl1_d3;
            ofl1_d5 <=  ofl1_d4;
            ofl3_d1 <=  ofl3;
            ofl3_d2 <=  ofl3_d1;
            ofl3_d3 <=  ofl3_d2;
            ofl3_d4 <=  ofl3_d3;
            ofl3_d5 <=  ofl3_d4;
            ofl3_d6 <=  ofl3_d5;
            ofl3_d7 <=  ofl3_d6;
            ufl2_d1 <=  ufl2;
            ufl2_d2 <=  ufl2_d1;
            ufl2_d3 <=  ufl2_d2;
            ufl2_d4 <=  ufl2_d3;
            ufl2_d5 <=  ufl2_d4;
            ufl2_d6 <=  ufl2_d5;
            ufl2_d7 <=  ufl2_d6;
            ufl3_d1 <=  ufl3;
            ufl3_d2 <=  ufl3_d1;
            ufl3_d3 <=  ufl3_d2;
            ufl3_d4 <=  ufl3_d3;
            ufl3_d5 <=  ufl3_d4;
         end if;
      end process;
   Xexn <= X(wE+wFIn+2 downto wE+wFIn+1);
   XSign <= X(wE+wFIn);
   XexpField <= X(wE+wFIn-1 downto wFIn);
   Xfrac <= unsigned(X(wFIn-1 downto 0));
   e0 <= conv_std_logic_vector(114, wE+2);  -- bias - (wF+g)
   shiftVal <= ("00" & XexpField_d1) - e0_d14; -- for a left shift
   -- underflow when input is shifted to zero (shiftval<0), in which case exp = 1
   resultWillBeOne <= shiftVal(wE+1);
   --  mantissa with implicit bit
   mXu <= "1" & Xfrac;
   -- Partial overflow detection
   maxShift <= conv_std_logic_vector(19, wE+1);  -- wE-2 + wF+g
   overflow0 <= not shiftVal_d1(wE+1) when shiftVal_d1(wE downto 0) > maxShift_d15 else '0';
   shiftValIn <= shiftVal(4 downto 0);
   mantissa_shift: LeftShifter22_by_max_19_Freq500_uid73
      port map ( clk  => clk,
                 S => shiftValIn,
                 X => std_logic_vector(mXu),
                 R => fixX0);
   ufixX <=  unsigned(fixX0(40 downto 21)) when resultWillBeOne_d1='0' else "00000000000000000000";
   exp_helper: Exp_8_10_Freq500_uid75
      port map ( clk  => clk,
                 XSign => XSign,
                 ufixX_i => std_logic_vector(ufixX),
                 K => K,
                 expY => expY);
   needNoNorm <= expY(13);
   -- Rounding: all this should consume one row of LUTs
   preRoundBiasSig <= conv_std_logic_vector(127, wE+2)  & expY(12 downto 3) when needNoNorm = '1'
      else conv_std_logic_vector(126, wE+2)  & expY(11 downto 2) ;
   roundBit <= expY(2)  when needNoNorm = '1'    else expY(1) ;
   roundNormAddend <= K_d2(8) & K_d2 & (9 downto 1 => '0') & roundBit;
   roundedExpSigOperandAdder: IntAdder_20_Freq500_uid121
      port map ( clk  => clk,
                 Cin => '0',
                 X => preRoundBiasSig,
                 Y => roundNormAddend,
                 R => roundedExpSigRes);
   roundedExpSig <= roundedExpSigRes when Xexn_d7="01" else  "000" & (wE-2 downto 0 => '1') & (wF-1 downto 0 => '0');
   ofl1 <= not XSign_d2 and overflow0 and (not Xexn_d2(1) and Xexn_d2(0)); -- input positive, normal,  very large
   ofl2 <= not XSign_d7 and (roundedExpSig(wE+wF) and not roundedExpSig(wE+wF+1)) and (not Xexn_d7(1) and Xexn_d7(0)); -- input positive, normal, overflowed
   ofl3 <= not XSign and Xexn(1) and not Xexn(0);  -- input was -infty
   ofl <= ofl1_d5 or ofl2 or ofl3_d7;
   ufl1 <= (roundedExpSig(wE+wF) and roundedExpSig(wE+wF+1))  and (not Xexn_d7(1) and Xexn_d7(0)); -- input normal
   ufl2 <= XSign and Xexn(1) and not Xexn(0);  -- input was -infty
   ufl3 <= XSign_d2 and overflow0  and (not Xexn_d2(1) and Xexn_d2(0)); -- input negative, normal,  very large
   ufl <= ufl1 or ufl2_d7 or ufl3_d5;
   Rexn <= "11" when Xexn_d7 = "11"
      else "10" when ofl='1'
      else "00" when ufl='1'
      else "01";
   R <= Rexn & '0' & roundedExpSig(17 downto 0);
end architecture;

--------------------------------------------------------------------------------
--                                 top_module
--                         (FPPow_8_10_Freq500_uid2)
-- VHDL generated for DummyFPGA @ 500MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: F. de Dinechin, C. Klein  (2008)
--------------------------------------------------------------------------------
-- Pipeline depth: 21 cycles
-- Clock period (ns): 2
-- Target frequency (MHz): 500
-- Input signals: X Y
-- Output signals: R
--  approx. input signal timings: X: (c0, 0.000000ns)Y: (c0, 0.000000ns)
--  approx. output signal timings: R: (c21, 1.539231ns)

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity top_module is
    port (clk : in std_logic;
          X : in  std_logic_vector(8+10+2 downto 0);
          Y : in  std_logic_vector(8+10+2 downto 0);
          R : out  std_logic_vector(8+10+2 downto 0)   );
end entity;

architecture arch of top_module is
   component IntAdder_19_Freq500_uid5 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(18 downto 0);
             Y : in  std_logic_vector(18 downto 0);
             Cin : in  std_logic;
             R : out  std_logic_vector(18 downto 0)   );
   end component;

   component LZC_10_Freq500_uid7 is
      port ( clk : in std_logic;
             I : in  std_logic_vector(9 downto 0);
             O : out  std_logic_vector(3 downto 0)   );
   end component;

   component FPLogIterative_8_20_0_500_Freq500_uid9 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(8+20+2 downto 0);
             R : out  std_logic_vector(8+20+2 downto 0)   );
   end component;

   component FPMult_8_20_uid62_Freq500_uid63 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(8+20+2 downto 0);
             Y : in  std_logic_vector(8+10+2 downto 0);
             R : out  std_logic_vector(8+21+2 downto 0)   );
   end component;

   component FPExp_8_10_Freq500_uid71 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(8+21+2 downto 0);
             R : out  std_logic_vector(8+10+2 downto 0)   );
   end component;

signal flagsX :  std_logic_vector(1 downto 0);
   -- timing of flagsX: (c0, 0.000000ns)
signal signX, signX_d1, signX_d2 :  std_logic;
   -- timing of signX: (c0, 0.000000ns)
signal expFieldX :  std_logic_vector(7 downto 0);
   -- timing of expFieldX: (c0, 0.000000ns)
signal fracX :  std_logic_vector(9 downto 0);
   -- timing of fracX: (c0, 0.000000ns)
signal flagsY :  std_logic_vector(1 downto 0);
   -- timing of flagsY: (c0, 0.000000ns)
signal signY, signY_d1, signY_d2, signY_d3 :  std_logic;
   -- timing of signY: (c0, 0.000000ns)
signal expFieldY :  std_logic_vector(7 downto 0);
   -- timing of expFieldY: (c0, 0.000000ns)
signal fracY :  std_logic_vector(9 downto 0);
   -- timing of fracY: (c0, 0.000000ns)
signal zeroX, zeroX_d1, zeroX_d2, zeroX_d3 :  std_logic;
   -- timing of zeroX: (c0, 0.550000ns)
signal zeroY, zeroY_d1, zeroY_d2 :  std_logic;
   -- timing of zeroY: (c0, 0.550000ns)
signal normalX, normalX_d1, normalX_d2 :  std_logic;
   -- timing of normalX: (c0, 0.550000ns)
signal normalY, normalY_d1, normalY_d2, normalY_d3 :  std_logic;
   -- timing of normalY: (c0, 0.550000ns)
signal infX, infX_d1, infX_d2, infX_d3 :  std_logic;
   -- timing of infX: (c0, 0.550000ns)
signal infY, infY_d1, infY_d2, infY_d3 :  std_logic;
   -- timing of infY: (c0, 0.550000ns)
signal s_nan_in, s_nan_in_d1, s_nan_in_d2 :  std_logic;
   -- timing of s_nan_in: (c0, 0.550000ns)
signal OneExpFrac :  std_logic_vector(17 downto 0);
   -- timing of OneExpFrac: (c0, 0.000000ns)
signal ExpFracX :  std_logic_vector(18 downto 0);
   -- timing of ExpFracX: (c0, 0.000000ns)
signal OneExpFracCompl :  std_logic_vector(18 downto 0);
   -- timing of OneExpFracCompl: (c0, 0.000000ns)
signal cmpXOneRes :  std_logic_vector(18 downto 0);
   -- timing of cmpXOneRes: (c0, 1.180000ns)
signal XisOneAndNormal :  std_logic;
   -- timing of XisOneAndNormal: (c0, 0.550000ns)
signal absXgtOneAndNormal, absXgtOneAndNormal_d1, absXgtOneAndNormal_d2, absXgtOneAndNormal_d3 :  std_logic;
   -- timing of absXgtOneAndNormal: (c0, 1.730000ns)
signal absXltOneAndNormal, absXltOneAndNormal_d1, absXltOneAndNormal_d2, absXltOneAndNormal_d3 :  std_logic;
   -- timing of absXltOneAndNormal: (c0, 1.730000ns)
signal fracYreverted :  std_logic_vector(9 downto 0);
   -- timing of fracYreverted: (c0, 0.000000ns)
signal Z_rightY, Z_rightY_d1 :  std_logic_vector(3 downto 0);
   -- timing of Z_rightY: (c1, 0.980000ns)
signal WeightLSBYpre, WeightLSBYpre_d1, WeightLSBYpre_d2 :  std_logic_vector(8 downto 0);
   -- timing of WeightLSBYpre: (c0, 1.080000ns)
signal WeightLSBY :  std_logic_vector(8 downto 0);
   -- timing of WeightLSBY: (c2, 0.260000ns)
signal oddIntY, oddIntY_d1 :  std_logic;
   -- timing of oddIntY: (c2, 0.810000ns)
signal evenIntY, evenIntY_d1 :  std_logic;
   -- timing of evenIntY: (c2, 1.360000ns)
signal notIntNormalY :  std_logic;
   -- timing of notIntNormalY: (c2, 0.810000ns)
signal RisInfSpecialCase, RisInfSpecialCase_d1, RisInfSpecialCase_d2, RisInfSpecialCase_d3, RisInfSpecialCase_d4, RisInfSpecialCase_d5, RisInfSpecialCase_d6, RisInfSpecialCase_d7, RisInfSpecialCase_d8, RisInfSpecialCase_d9, RisInfSpecialCase_d10, RisInfSpecialCase_d11, RisInfSpecialCase_d12, RisInfSpecialCase_d13, RisInfSpecialCase_d14, RisInfSpecialCase_d15, RisInfSpecialCase_d16, RisInfSpecialCase_d17, RisInfSpecialCase_d18 :  std_logic;
   -- timing of RisInfSpecialCase: (c3, 0.110000ns)
signal RisZeroSpecialCase, RisZeroSpecialCase_d1, RisZeroSpecialCase_d2, RisZeroSpecialCase_d3, RisZeroSpecialCase_d4, RisZeroSpecialCase_d5, RisZeroSpecialCase_d6, RisZeroSpecialCase_d7, RisZeroSpecialCase_d8, RisZeroSpecialCase_d9, RisZeroSpecialCase_d10, RisZeroSpecialCase_d11, RisZeroSpecialCase_d12, RisZeroSpecialCase_d13, RisZeroSpecialCase_d14, RisZeroSpecialCase_d15, RisZeroSpecialCase_d16, RisZeroSpecialCase_d17, RisZeroSpecialCase_d18 :  std_logic;
   -- timing of RisZeroSpecialCase: (c3, 0.110000ns)
signal RisOne, RisOne_d1, RisOne_d2, RisOne_d3, RisOne_d4, RisOne_d5, RisOne_d6, RisOne_d7, RisOne_d8, RisOne_d9, RisOne_d10, RisOne_d11, RisOne_d12, RisOne_d13, RisOne_d14, RisOne_d15, RisOne_d16, RisOne_d17, RisOne_d18, RisOne_d19, RisOne_d20, RisOne_d21 :  std_logic;
   -- timing of RisOne: (c0, 1.100000ns)
signal RisNaN, RisNaN_d1, RisNaN_d2, RisNaN_d3, RisNaN_d4, RisNaN_d5, RisNaN_d6, RisNaN_d7, RisNaN_d8, RisNaN_d9, RisNaN_d10, RisNaN_d11, RisNaN_d12, RisNaN_d13, RisNaN_d14, RisNaN_d15, RisNaN_d16, RisNaN_d17, RisNaN_d18, RisNaN_d19 :  std_logic;
   -- timing of RisNaN: (c2, 0.810000ns)
signal signR, signR_d1, signR_d2, signR_d3, signR_d4, signR_d5, signR_d6, signR_d7, signR_d8, signR_d9, signR_d10, signR_d11, signR_d12, signR_d13, signR_d14, signR_d15, signR_d16, signR_d17, signR_d18, signR_d19 :  std_logic;
   -- timing of signR: (c2, 0.810000ns)
signal logIn :  std_logic_vector(30 downto 0);
   -- timing of logIn: (c0, 0.000000ns)
signal lnX :  std_logic_vector(8+20+2 downto 0);
   -- timing of lnX: (c11, 1.735385ns)
signal P :  std_logic_vector(8+21+2 downto 0);
   -- timing of P: (c13, 1.615385ns)
signal E, E_d1 :  std_logic_vector(8+10+2 downto 0);
   -- timing of E: (c20, 1.689231ns)
signal flagsE, flagsE_d1 :  std_logic_vector(1 downto 0);
   -- timing of flagsE: (c20, 1.689231ns)
signal RisZeroFromExp :  std_logic;
   -- timing of RisZeroFromExp: (c21, 0.439231ns)
signal RisZero :  std_logic;
   -- timing of RisZero: (c21, 0.989231ns)
signal RisInfFromExp :  std_logic;
   -- timing of RisInfFromExp: (c21, 0.439231ns)
signal RisInf :  std_logic;
   -- timing of RisInf: (c21, 0.989231ns)
signal flagR :  std_logic_vector(1 downto 0);
   -- timing of flagR: (c21, 1.539231ns)
signal R_expfrac :  std_logic_vector(17 downto 0);
   -- timing of R_expfrac: (c21, 0.439231ns)
constant wE: positive := 8;
constant wF: positive := 10;
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            signX_d1 <=  signX;
            signX_d2 <=  signX_d1;
            signY_d1 <=  signY;
            signY_d2 <=  signY_d1;
            signY_d3 <=  signY_d2;
            zeroX_d1 <=  zeroX;
            zeroX_d2 <=  zeroX_d1;
            zeroX_d3 <=  zeroX_d2;
            zeroY_d1 <=  zeroY;
            zeroY_d2 <=  zeroY_d1;
            normalX_d1 <=  normalX;
            normalX_d2 <=  normalX_d1;
            normalY_d1 <=  normalY;
            normalY_d2 <=  normalY_d1;
            normalY_d3 <=  normalY_d2;
            infX_d1 <=  infX;
            infX_d2 <=  infX_d1;
            infX_d3 <=  infX_d2;
            infY_d1 <=  infY;
            infY_d2 <=  infY_d1;
            infY_d3 <=  infY_d2;
            s_nan_in_d1 <=  s_nan_in;
            s_nan_in_d2 <=  s_nan_in_d1;
            absXgtOneAndNormal_d1 <=  absXgtOneAndNormal;
            absXgtOneAndNormal_d2 <=  absXgtOneAndNormal_d1;
            absXgtOneAndNormal_d3 <=  absXgtOneAndNormal_d2;
            absXltOneAndNormal_d1 <=  absXltOneAndNormal;
            absXltOneAndNormal_d2 <=  absXltOneAndNormal_d1;
            absXltOneAndNormal_d3 <=  absXltOneAndNormal_d2;
            Z_rightY_d1 <=  Z_rightY;
            WeightLSBYpre_d1 <=  WeightLSBYpre;
            WeightLSBYpre_d2 <=  WeightLSBYpre_d1;
            oddIntY_d1 <=  oddIntY;
            evenIntY_d1 <=  evenIntY;
            RisInfSpecialCase_d1 <=  RisInfSpecialCase;
            RisInfSpecialCase_d2 <=  RisInfSpecialCase_d1;
            RisInfSpecialCase_d3 <=  RisInfSpecialCase_d2;
            RisInfSpecialCase_d4 <=  RisInfSpecialCase_d3;
            RisInfSpecialCase_d5 <=  RisInfSpecialCase_d4;
            RisInfSpecialCase_d6 <=  RisInfSpecialCase_d5;
            RisInfSpecialCase_d7 <=  RisInfSpecialCase_d6;
            RisInfSpecialCase_d8 <=  RisInfSpecialCase_d7;
            RisInfSpecialCase_d9 <=  RisInfSpecialCase_d8;
            RisInfSpecialCase_d10 <=  RisInfSpecialCase_d9;
            RisInfSpecialCase_d11 <=  RisInfSpecialCase_d10;
            RisInfSpecialCase_d12 <=  RisInfSpecialCase_d11;
            RisInfSpecialCase_d13 <=  RisInfSpecialCase_d12;
            RisInfSpecialCase_d14 <=  RisInfSpecialCase_d13;
            RisInfSpecialCase_d15 <=  RisInfSpecialCase_d14;
            RisInfSpecialCase_d16 <=  RisInfSpecialCase_d15;
            RisInfSpecialCase_d17 <=  RisInfSpecialCase_d16;
            RisInfSpecialCase_d18 <=  RisInfSpecialCase_d17;
            RisZeroSpecialCase_d1 <=  RisZeroSpecialCase;
            RisZeroSpecialCase_d2 <=  RisZeroSpecialCase_d1;
            RisZeroSpecialCase_d3 <=  RisZeroSpecialCase_d2;
            RisZeroSpecialCase_d4 <=  RisZeroSpecialCase_d3;
            RisZeroSpecialCase_d5 <=  RisZeroSpecialCase_d4;
            RisZeroSpecialCase_d6 <=  RisZeroSpecialCase_d5;
            RisZeroSpecialCase_d7 <=  RisZeroSpecialCase_d6;
            RisZeroSpecialCase_d8 <=  RisZeroSpecialCase_d7;
            RisZeroSpecialCase_d9 <=  RisZeroSpecialCase_d8;
            RisZeroSpecialCase_d10 <=  RisZeroSpecialCase_d9;
            RisZeroSpecialCase_d11 <=  RisZeroSpecialCase_d10;
            RisZeroSpecialCase_d12 <=  RisZeroSpecialCase_d11;
            RisZeroSpecialCase_d13 <=  RisZeroSpecialCase_d12;
            RisZeroSpecialCase_d14 <=  RisZeroSpecialCase_d13;
            RisZeroSpecialCase_d15 <=  RisZeroSpecialCase_d14;
            RisZeroSpecialCase_d16 <=  RisZeroSpecialCase_d15;
            RisZeroSpecialCase_d17 <=  RisZeroSpecialCase_d16;
            RisZeroSpecialCase_d18 <=  RisZeroSpecialCase_d17;
            RisOne_d1 <=  RisOne;
            RisOne_d2 <=  RisOne_d1;
            RisOne_d3 <=  RisOne_d2;
            RisOne_d4 <=  RisOne_d3;
            RisOne_d5 <=  RisOne_d4;
            RisOne_d6 <=  RisOne_d5;
            RisOne_d7 <=  RisOne_d6;
            RisOne_d8 <=  RisOne_d7;
            RisOne_d9 <=  RisOne_d8;
            RisOne_d10 <=  RisOne_d9;
            RisOne_d11 <=  RisOne_d10;
            RisOne_d12 <=  RisOne_d11;
            RisOne_d13 <=  RisOne_d12;
            RisOne_d14 <=  RisOne_d13;
            RisOne_d15 <=  RisOne_d14;
            RisOne_d16 <=  RisOne_d15;
            RisOne_d17 <=  RisOne_d16;
            RisOne_d18 <=  RisOne_d17;
            RisOne_d19 <=  RisOne_d18;
            RisOne_d20 <=  RisOne_d19;
            RisOne_d21 <=  RisOne_d20;
            RisNaN_d1 <=  RisNaN;
            RisNaN_d2 <=  RisNaN_d1;
            RisNaN_d3 <=  RisNaN_d2;
            RisNaN_d4 <=  RisNaN_d3;
            RisNaN_d5 <=  RisNaN_d4;
            RisNaN_d6 <=  RisNaN_d5;
            RisNaN_d7 <=  RisNaN_d6;
            RisNaN_d8 <=  RisNaN_d7;
            RisNaN_d9 <=  RisNaN_d8;
            RisNaN_d10 <=  RisNaN_d9;
            RisNaN_d11 <=  RisNaN_d10;
            RisNaN_d12 <=  RisNaN_d11;
            RisNaN_d13 <=  RisNaN_d12;
            RisNaN_d14 <=  RisNaN_d13;
            RisNaN_d15 <=  RisNaN_d14;
            RisNaN_d16 <=  RisNaN_d15;
            RisNaN_d17 <=  RisNaN_d16;
            RisNaN_d18 <=  RisNaN_d17;
            RisNaN_d19 <=  RisNaN_d18;
            signR_d1 <=  signR;
            signR_d2 <=  signR_d1;
            signR_d3 <=  signR_d2;
            signR_d4 <=  signR_d3;
            signR_d5 <=  signR_d4;
            signR_d6 <=  signR_d5;
            signR_d7 <=  signR_d6;
            signR_d8 <=  signR_d7;
            signR_d9 <=  signR_d8;
            signR_d10 <=  signR_d9;
            signR_d11 <=  signR_d10;
            signR_d12 <=  signR_d11;
            signR_d13 <=  signR_d12;
            signR_d14 <=  signR_d13;
            signR_d15 <=  signR_d14;
            signR_d16 <=  signR_d15;
            signR_d17 <=  signR_d16;
            signR_d18 <=  signR_d17;
            signR_d19 <=  signR_d18;
            E_d1 <=  E;
            flagsE_d1 <=  flagsE;
         end if;
      end process;
   flagsX <= X(wE+wF+2 downto wE+wF+1);
   signX <= X(wE+wF);
   expFieldX <= X(wE+wF-1 downto wF);
   fracX <= X(wF-1 downto 0);
   flagsY <= Y(wE+wF+2 downto wE+wF+1);
   signY <= Y(wE+wF);
   expFieldY <= Y(wE+wF-1 downto wF);
   fracY <= Y(wF-1 downto 0);
-- Inputs analysis  --
-- zero inputs--
   zeroX <= '1' when flagsX="00" else '0';
   zeroY <= '1' when flagsY="00" else '0';
-- normal inputs--
   normalX <= '1' when flagsX="01" else '0';
   normalY <= '1' when flagsY="01" else '0';
-- inf input --
   infX <= '1' when flagsX="10" else '0';
   infY <= '1' when flagsY="10" else '0';
-- NaN inputs  --
   s_nan_in <= '1' when flagsX="11" or flagsY="11" else '0';
-- Comparison of X to 1   --
   OneExpFrac <=  "0" & (6 downto 0 => '1') & (9 downto 0 => '0');
   ExpFracX<= "0" & expFieldX & fracX;
   OneExpFracCompl<=  "1" & (not OneExpFrac);
   cmpXOne: IntAdder_19_Freq500_uid5
      port map ( clk  => clk,
                 Cin => '1',
                 X => ExpFracX,
                 Y => OneExpFracCompl,
                 R => cmpXOneRes);
   XisOneAndNormal <= '1' when X = ("010" & OneExpFrac) else '0';
   absXgtOneAndNormal <= normalX and (not XisOneAndNormal) and (not cmpXOneRes(18));
   absXltOneAndNormal <= normalX and cmpXOneRes(18);
   fracYreverted <= fracY(0)&fracY(1)&fracY(2)&fracY(3)&fracY(4)&fracY(5)&fracY(6)&fracY(7)&fracY(8)&fracY(9);
   FPPow_8_10_Freq500_uid2right1counter: LZC_10_Freq500_uid7
      port map ( clk  => clk,
                 I => fracYreverted,
                 O => Z_rightY);
-- compute the weight of the less significant one of the mantissa
   WeightLSBYpre <= ('0' & expFieldY)- CONV_STD_LOGIC_VECTOR(137,9);
   WeightLSBY <= WeightLSBYpre_d2 + Z_rightY_d1;
   oddIntY <= normalY_d2 when WeightLSBY = CONV_STD_LOGIC_VECTOR(0, 9) else '0'; -- LSB has null weight
   evenIntY <= normalY_d2 when WeightLSBY(wE)='0' and oddIntY='0' else '0'; --LSB has strictly positive weight 
   notIntNormalY <= normalY_d2 when WeightLSBY(wE)='1' else '0'; -- LSB has negative weight

-- Pow Exceptions  --
   RisInfSpecialCase  <= 
         (zeroX_d3  and  (oddIntY_d1 or evenIntY_d1)  and signY_d3)  -- (+/- 0) ^ (negative int y)
      or (zeroX_d3 and infY_d3 and signY_d3)                      -- (+/- 0) ^ (-inf)
      or (absXgtOneAndNormal_d3   and  infY_d3  and not signY_d3) -- (|x|>1) ^ (+inf)
      or (absXltOneAndNormal_d3   and  infY_d3  and signY_d3)     -- (|x|<1) ^ (-inf)
      or (infX_d3 and  normalY_d3  and not signY_d3) ;            -- (inf) ^ (y>0)
   RisZeroSpecialCase <= 
         (zeroX_d3 and  (oddIntY_d1 or evenIntY_d1)  and not signY_d3)  -- (+/- 0) ^ (positive int y)
      or (zeroX_d3 and  infY_d3  and not signY_d3)                   -- (+/- 0) ^ (+inf)
      or (absXltOneAndNormal_d3   and  infY_d3  and not signY_d3)    -- (|x|<1) ^ (+inf)
      or (absXgtOneAndNormal_d3   and  infY_d3  and signY_d3)        -- (|x|>1) ^ (-inf)
      or (infX_d3 and  normalY_d3  and signY_d3) ;                   -- (inf) ^ (y<0)
   RisOne <= 
         zeroY                                          -- x^0 = 1 without exception
      or (XisOneAndNormal and signX and infY)           -- (-1) ^ (-/-inf)
      or (XisOneAndNormal  and not signX);              -- (+1) ^ (whatever)
   RisNaN <= (s_nan_in_d2 and not zeroY_d2) or (normalX_d2 and signX_d2 and notIntNormalY);
   signR <= signX_d2 and (oddIntY);
   logIn <= flagsX & "0" & expFieldX & fracX & (9 downto 0 => '0') ;
   FPPow_8_10_Freq500_uid2log: FPLogIterative_8_20_0_500_Freq500_uid9
      port map ( clk  => clk,
                 X => logIn,
                 R => lnX);
   FPPow_8_10_Freq500_uid2mult: FPMult_8_20_uid62_Freq500_uid63
      port map ( clk  => clk,
                 X => lnX,
                 Y => Y,
                 R => P);
   FPPow_8_10_Freq500_uid2exp: FPExp_8_10_Freq500_uid71
      port map ( clk  => clk,
                 X => P,
                 R => E);
   flagsE <= E(wE+wF+2 downto wE+wF+1);
   RisZeroFromExp <= '1' when flagsE_d1="00" else '0';
   RisZero <= RisZeroSpecialCase_d18 or RisZeroFromExp;
   RisInfFromExp  <= '1' when flagsE_d1="10" else '0';
   RisInf  <= RisInfSpecialCase_d18 or RisInfFromExp;
   flagR <= 
           "11" when RisNaN_d19='1'
      else "00" when RisZero='1'
      else "10" when RisInf='1'
      else "01";
   R_expfrac <= CONV_STD_LOGIC_VECTOR(127,8) &  CONV_STD_LOGIC_VECTOR(0, 10) when RisOne_d21='1'
       else E_d1(17 downto 0);
   R <= flagR & signR_d19 & R_expfrac;
end architecture;

--------------------------------------------------------------------------------
--                    TestBench_top_module_Freq500_uid123
-- VHDL generated for DummyFPGA @ 500MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Cristian Klein, Nicolas Brunie (2007-2010)
--------------------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity TestBench_top_module_Freq500_uid123 is
end entity;

architecture behavorial of TestBench_top_module_Freq500_uid123 is
   component top_module is
      port ( clk : in std_logic;
             X : in  std_logic_vector(8+10+2 downto 0);
             Y : in  std_logic_vector(8+10+2 downto 0);
             R : out  std_logic_vector(8+10+2 downto 0)   );
   end component;
signal X :  std_logic_vector(20 downto 0);
   -- timing of X: (c0, 0.000000ns)
signal Y :  std_logic_vector(20 downto 0);
   -- timing of Y: (c0, 0.000000ns)
signal R :  std_logic_vector(20 downto 0);
   -- timing of R: (c21, 0.000000ns)
signal clk :  std_logic;
   -- timing of clk: (c0, 0.000000ns)
signal rst :  std_logic;
   -- timing of rst: (c0, 0.000000ns)

 -- converts std_logic into a character
   function chr(sl: std_logic) return character is
      variable c: character;
   begin
      case sl is
         when 'U' => c:= 'U';
         when 'X' => c:= 'X';
         when '0' => c:= '0';
         when '1' => c:= '1';
         when 'Z' => c:= 'Z';
         when 'W' => c:= 'W';
         when 'L' => c:= 'L';
         when 'H' => c:= 'H';
         when '-' => c:= '-';
      end case;
      return c;
   end chr;

   -- converts bit to std_logic (1 to 1)
   function to_stdlogic(b : bit) return std_logic is
       variable sl : std_logic;
   begin
      case b is 
         when '0' => sl := '0';
         when '1' => sl := '1';
      end case;
      return sl;
   end to_stdlogic;

   -- converts std_logic into a string (1 to 1)
   function str(sl: std_logic) return string is
    variable s: string(1 to 1);
    begin
      s(1) := chr(sl);
      return s;
   end str;

   -- converts std_logic_vector into a string (binary base)
   -- (this also takes care of the fact that the range of
   --  a string is natural while a std_logic_vector may
   --  have an integer range)
   function str(slv: std_logic_vector) return string is
      variable result : string (1 to slv'length);
      variable r : integer;
   begin
      r := 1;
      for i in slv'range loop
         result(r) := chr(slv(i));
         r := r + 1;
      end loop;
      return result;
   end str;

   -- FP compare function (found vs. real)
   function fp_equal(a : std_logic_vector; b : std_logic_vector) return boolean is
   begin
      if b(b'high downto b'high-1) = "01" then
         return a = b;
      elsif b(b'high downto b'high-1) = "11" then
         return (a(a'high downto a'high-1)=b(b'high downto b'high-1));
      else
         return a(a'high downto a'high-2) = b(b'high downto b'high-2);
      end if;
   end;

   function fp_inf_or_equal(a : std_logic_vector; b : std_logic_vector) return boolean is
   begin
      if (b(b'high downto b'high-1) = "11") or (a(a'high downto a'high-1) = "11")  then
         return false; -- NaN always compare false
      else return true; -- TODO
      end if;
   end;

   -- FP subtypes for casting
   subtype fp21 is std_logic_vector(20 downto 0);
   function testLine(testCounter:integer; expectedOutputS: string(1 to 10000); expectedOutputSize: integer; R:  std_logic_vector(8+10+2 downto 0)) return boolean is
      variable expectedOutput: line;
      variable possibilityNumber : integer;
      variable testSuccess: boolean;
      variable errorMessage: string(1 to 10000);
      variable testSuccess_R: boolean;
      variable expected_R: bit_vector (20 downto 0); -- for list of values
      variable inf_R: bit_vector (20 downto 0); -- for intervals
      variable sup_R: bit_vector (20 downto 0); -- for intervals
   begin
      write(expectedOutput, expectedOutputS);
      read(expectedOutput, possibilityNumber); -- for R
      if possibilityNumber = 0 then
         -- TODO define what it means to have 0 possible output. Currently it means a test fails...
      end if;
      if possibilityNumber > 0 then -- a list of values
      testSuccess_R := false;
         for i in 1 to possibilityNumber loop
            read(expectedOutput, expected_R);
            if fp_equal(R, to_stdlogicvector(expected_R)) then
               testSuccess_R := true;
            end if;
            end loop;
      end if;
      if possibilityNumber < 0  then -- an interval
         read(expectedOutput, inf_R);
         read(expectedOutput, sup_R);
         if possibilityNumber =-1  then -- an unsigned interval
            testSuccess_R := (R >= to_stdlogicvector(inf_R)) and (R <= to_stdlogicvector(sup_R));
         elsif possibilityNumber =-2  then -- a signed interval
            testSuccess_R := (signed(R) >= signed(to_stdlogicvector(inf_R))) and (signed(R) <= signed(to_stdlogicvector(sup_R)));
         elsif possibilityNumber =-4  then -- a floating-point interval
            testSuccess_R := fp_inf_or_equal(to_stdlogicvector(inf_R), R) and fp_inf_or_equal(R, to_stdlogicvector(sup_R));
         end if;
      end if;
      if testSuccess_R = false then
         report("Test #" & integer'image(testCounter) & ", incorrect output for R: " & lf & " expected values: " & expectedOutputS(1 to expectedOutputSize) & lf  & "          result:    " & str(R) ) severity error;
      end if;
      
      testSuccess := true and testSuccess_R;
      return testSuccess;
   end testLine;

begin
   -- Ticking clock signal
   process
   begin
      clk <= '0';
      wait for 5 ns;
      clk <= '1';
      wait for 5 ns;
   end process;

   test: top_module
      port map ( clk  => clk,
                 X => X,
                 Y => Y,
                 R => R);
   -- Process that sets the inputs  (read from a file) 
   process
      variable input, expectedOutput : line; 
      variable tmpChar : character;
      file inputsFile : text is "test.input"; 
      variable V_X : bit_vector(20 downto 0);
      variable V_Y : bit_vector(20 downto 0);
      variable V_R : bit_vector(20 downto 0);
   begin
      -- Send reset
      rst <= '1';
      wait for 10 ns;
      rst <= '0';
      readline(inputsFile, input); -- skip the first line of advertising
      while not endfile(inputsFile) loop
         readline(inputsFile, input); -- skip the comment line
         readline(inputsFile, input);
         readline(inputsFile, expectedOutput); -- comment line, unused in this process
         readline(inputsFile, expectedOutput); -- unused in this process
         read(input ,V_X);
         read(input,tmpChar);
         X <= to_stdlogicvector(V_X);
         read(input ,V_Y);
         read(input,tmpChar);
         Y <= to_stdlogicvector(V_Y);
         wait for 10 ns;
      end loop;
         wait for 310 ns; -- wait for pipeline to flush (and some more)
   end process;

    -- Process that verifies the corresponding output
   process
      file inputsFile : text is "test.input"; 
      variable input, expectedOutput : line; 
      variable testCounter : integer := 1;
      variable errorCounter : integer := 0;
      variable expectedOutputString : string(1 to 10000);
      variable testSuccess: boolean;
   begin
      wait for 12 ns; -- wait for reset 
      wait for 210 ns; -- wait for pipeline to flush
      readline(inputsFile, input); -- skip the first line of advertising
      while not endfile(inputsFile) loop
         readline(inputsFile, input); -- input comment, unused
         readline(inputsFile, input); -- input line, unused
         readline(inputsFile, expectedOutput); -- comment line, unused in this process
         readline(inputsFile, expectedOutput);
         expectedOutputString := expectedOutput.all & (expectedOutput'Length+1 to 10000 => ' ');
         testSuccess := testLine(testCounter, expectedOutputString, expectedOutput'Length, R);
         if not testSuccess then 
               errorCounter := errorCounter + 1; -- incrementing global error counter
         end if;
            testCounter := testCounter + 1; -- incrementing global error counter
         wait for 10 ns;
      end loop;
      report integer'image(errorCounter) & " error(s) encoutered." severity note;
      report "End of simulation after " & integer'image(testCounter-1) & " tests" severity note;
   end process;

end architecture;

