module intadder_18_freq500_uid99
  (input  clk,
   input  [17:0] x,
   input  [17:0] y,
   input  cin,
   output [17:0] r);
  wire [17:0] rtmp;
  wire [17:0] x_d1;
  wire [17:0] y_d1;
  wire cin_d1;
  wire cin_d2;
  wire cin_d3;
  wire cin_d4;
  wire cin_d5;
  wire cin_d6;
  wire cin_d7;
  wire cin_d8;
  wire cin_d9;
  wire cin_d10;
  wire cin_d11;
  wire cin_d12;
  wire cin_d13;
  wire cin_d14;
  wire cin_d15;
  wire cin_d16;
  wire cin_d17;
  wire [17:0] n6551;
  wire [17:0] n6552;
  wire [17:0] n6553;
  reg [17:0] n6554;
  reg [17:0] n6555;
  reg n6556;
  reg n6557;
  reg n6558;
  reg n6559;
  reg n6560;
  reg n6561;
  reg n6562;
  reg n6563;
  reg n6564;
  reg n6565;
  reg n6566;
  reg n6567;
  reg n6568;
  reg n6569;
  reg n6570;
  reg n6571;
  reg n6572;
  assign r = rtmp; //(module output)
  /* fppowbf16.vhdl:4299:8  */
  assign rtmp = n6553; // (signal)
  /* fppowbf16.vhdl:4301:8  */
  assign x_d1 = n6554; // (signal)
  /* fppowbf16.vhdl:4303:8  */
  assign y_d1 = n6555; // (signal)
  /* fppowbf16.vhdl:4305:8  */
  assign cin_d1 = n6556; // (signal)
  /* fppowbf16.vhdl:4305:16  */
  assign cin_d2 = n6557; // (signal)
  /* fppowbf16.vhdl:4305:24  */
  assign cin_d3 = n6558; // (signal)
  /* fppowbf16.vhdl:4305:32  */
  assign cin_d4 = n6559; // (signal)
  /* fppowbf16.vhdl:4305:40  */
  assign cin_d5 = n6560; // (signal)
  /* fppowbf16.vhdl:4305:48  */
  assign cin_d6 = n6561; // (signal)
  /* fppowbf16.vhdl:4305:56  */
  assign cin_d7 = n6562; // (signal)
  /* fppowbf16.vhdl:4305:64  */
  assign cin_d8 = n6563; // (signal)
  /* fppowbf16.vhdl:4305:72  */
  assign cin_d9 = n6564; // (signal)
  /* fppowbf16.vhdl:4305:80  */
  assign cin_d10 = n6565; // (signal)
  /* fppowbf16.vhdl:4305:89  */
  assign cin_d11 = n6566; // (signal)
  /* fppowbf16.vhdl:4305:98  */
  assign cin_d12 = n6567; // (signal)
  /* fppowbf16.vhdl:4305:107  */
  assign cin_d13 = n6568; // (signal)
  /* fppowbf16.vhdl:4305:116  */
  assign cin_d14 = n6569; // (signal)
  /* fppowbf16.vhdl:4305:125  */
  assign cin_d15 = n6570; // (signal)
  /* fppowbf16.vhdl:4305:134  */
  assign cin_d16 = n6571; // (signal)
  /* fppowbf16.vhdl:4305:143  */
  assign cin_d17 = n6572; // (signal)
  /* fppowbf16.vhdl:4332:17  */
  assign n6551 = x_d1 + y_d1;
  /* fppowbf16.vhdl:4332:24  */
  assign n6552 = {17'b0, cin_d17};  //  uext
  /* fppowbf16.vhdl:4332:24  */
  assign n6553 = n6551 + n6552;
  /* fppowbf16.vhdl:4310:10  */
  always @(posedge clk)
    n6554 <= x;
  /* fppowbf16.vhdl:4310:10  */
  always @(posedge clk)
    n6555 <= y;
  /* fppowbf16.vhdl:4310:10  */
  always @(posedge clk)
    n6556 <= cin;
  /* fppowbf16.vhdl:4310:10  */
  always @(posedge clk)
    n6557 <= cin_d1;
  /* fppowbf16.vhdl:4310:10  */
  always @(posedge clk)
    n6558 <= cin_d2;
  /* fppowbf16.vhdl:4310:10  */
  always @(posedge clk)
    n6559 <= cin_d3;
  /* fppowbf16.vhdl:4310:10  */
  always @(posedge clk)
    n6560 <= cin_d4;
  /* fppowbf16.vhdl:4310:10  */
  always @(posedge clk)
    n6561 <= cin_d5;
  /* fppowbf16.vhdl:4310:10  */
  always @(posedge clk)
    n6562 <= cin_d6;
  /* fppowbf16.vhdl:4310:10  */
  always @(posedge clk)
    n6563 <= cin_d7;
  /* fppowbf16.vhdl:4310:10  */
  always @(posedge clk)
    n6564 <= cin_d8;
  /* fppowbf16.vhdl:4310:10  */
  always @(posedge clk)
    n6565 <= cin_d9;
  /* fppowbf16.vhdl:4310:10  */
  always @(posedge clk)
    n6566 <= cin_d10;
  /* fppowbf16.vhdl:4310:10  */
  always @(posedge clk)
    n6567 <= cin_d11;
  /* fppowbf16.vhdl:4310:10  */
  always @(posedge clk)
    n6568 <= cin_d12;
  /* fppowbf16.vhdl:4310:10  */
  always @(posedge clk)
    n6569 <= cin_d13;
  /* fppowbf16.vhdl:4310:10  */
  always @(posedge clk)
    n6570 <= cin_d14;
  /* fppowbf16.vhdl:4310:10  */
  always @(posedge clk)
    n6571 <= cin_d15;
  /* fppowbf16.vhdl:4310:10  */
  always @(posedge clk)
    n6572 <= cin_d16;
endmodule

module fixrealkcm_freq500_uid89_t1_freq500_uid95
  (input  [2:0] x,
   output [12:0] y);
  wire [12:0] y0;
  wire [12:0] y1;
  wire n6502;
  wire n6505;
  wire n6508;
  wire n6511;
  wire n6514;
  wire n6517;
  wire n6520;
  wire n6523;
  wire [7:0] n6525;
  reg [12:0] n6526;
  assign y = y1; //(module output)
  /* fppowbf16.vhdl:774:8  */
  assign y0 = n6526; // (signal)
  /* fppowbf16.vhdl:776:8  */
  assign y1 = y0; // (signal)
  /* fppowbf16.vhdl:780:23  */
  assign n6502 = x == 3'b000;
  /* fppowbf16.vhdl:781:23  */
  assign n6505 = x == 3'b001;
  /* fppowbf16.vhdl:782:23  */
  assign n6508 = x == 3'b010;
  /* fppowbf16.vhdl:783:23  */
  assign n6511 = x == 3'b011;
  /* fppowbf16.vhdl:784:23  */
  assign n6514 = x == 3'b100;
  /* fppowbf16.vhdl:785:23  */
  assign n6517 = x == 3'b101;
  /* fppowbf16.vhdl:786:23  */
  assign n6520 = x == 3'b110;
  /* fppowbf16.vhdl:787:23  */
  assign n6523 = x == 3'b111;
  assign n6525 = {n6523, n6520, n6517, n6514, n6511, n6508, n6505, n6502};
  /* fppowbf16.vhdl:779:4  */
  always @*
    case (n6525)
      8'b10000000: n6526 = 13'b1001101101000;
      8'b01000000: n6526 = 13'b1000010100011;
      8'b00100000: n6526 = 13'b0110111011101;
      8'b00010000: n6526 = 13'b0101100010111;
      8'b00001000: n6526 = 13'b0100001010001;
      8'b00000100: n6526 = 13'b0010110001100;
      8'b00000010: n6526 = 13'b0001011000110;
      8'b00000001: n6526 = 13'b0000000000000;
      default: n6526 = 13'bX;
    endcase
endmodule

module fixrealkcm_freq500_uid89_t0_freq500_uid92
  (input  [4:0] x,
   output [17:0] y);
  wire [17:0] y0;
  wire [17:0] y1;
  wire n6402;
  wire n6405;
  wire n6408;
  wire n6411;
  wire n6414;
  wire n6417;
  wire n6420;
  wire n6423;
  wire n6426;
  wire n6429;
  wire n6432;
  wire n6435;
  wire n6438;
  wire n6441;
  wire n6444;
  wire n6447;
  wire n6450;
  wire n6453;
  wire n6456;
  wire n6459;
  wire n6462;
  wire n6465;
  wire n6468;
  wire n6471;
  wire n6474;
  wire n6477;
  wire n6480;
  wire n6483;
  wire n6486;
  wire n6489;
  wire n6492;
  wire n6495;
  wire [31:0] n6497;
  reg [17:0] n6498;
  assign y = y1; //(module output)
  /* fppowbf16.vhdl:702:8  */
  assign y0 = n6498; // (signal)
  /* fppowbf16.vhdl:704:8  */
  assign y1 = y0; // (signal)
  /* fppowbf16.vhdl:708:28  */
  assign n6402 = x == 5'b00000;
  /* fppowbf16.vhdl:709:28  */
  assign n6405 = x == 5'b00001;
  /* fppowbf16.vhdl:710:28  */
  assign n6408 = x == 5'b00010;
  /* fppowbf16.vhdl:711:28  */
  assign n6411 = x == 5'b00011;
  /* fppowbf16.vhdl:712:28  */
  assign n6414 = x == 5'b00100;
  /* fppowbf16.vhdl:713:28  */
  assign n6417 = x == 5'b00101;
  /* fppowbf16.vhdl:714:28  */
  assign n6420 = x == 5'b00110;
  /* fppowbf16.vhdl:715:28  */
  assign n6423 = x == 5'b00111;
  /* fppowbf16.vhdl:716:28  */
  assign n6426 = x == 5'b01000;
  /* fppowbf16.vhdl:717:28  */
  assign n6429 = x == 5'b01001;
  /* fppowbf16.vhdl:718:28  */
  assign n6432 = x == 5'b01010;
  /* fppowbf16.vhdl:719:28  */
  assign n6435 = x == 5'b01011;
  /* fppowbf16.vhdl:720:28  */
  assign n6438 = x == 5'b01100;
  /* fppowbf16.vhdl:721:28  */
  assign n6441 = x == 5'b01101;
  /* fppowbf16.vhdl:722:28  */
  assign n6444 = x == 5'b01110;
  /* fppowbf16.vhdl:723:28  */
  assign n6447 = x == 5'b01111;
  /* fppowbf16.vhdl:724:28  */
  assign n6450 = x == 5'b10000;
  /* fppowbf16.vhdl:725:28  */
  assign n6453 = x == 5'b10001;
  /* fppowbf16.vhdl:726:28  */
  assign n6456 = x == 5'b10010;
  /* fppowbf16.vhdl:727:28  */
  assign n6459 = x == 5'b10011;
  /* fppowbf16.vhdl:728:28  */
  assign n6462 = x == 5'b10100;
  /* fppowbf16.vhdl:729:28  */
  assign n6465 = x == 5'b10101;
  /* fppowbf16.vhdl:730:28  */
  assign n6468 = x == 5'b10110;
  /* fppowbf16.vhdl:731:28  */
  assign n6471 = x == 5'b10111;
  /* fppowbf16.vhdl:732:28  */
  assign n6474 = x == 5'b11000;
  /* fppowbf16.vhdl:733:28  */
  assign n6477 = x == 5'b11001;
  /* fppowbf16.vhdl:734:28  */
  assign n6480 = x == 5'b11010;
  /* fppowbf16.vhdl:735:28  */
  assign n6483 = x == 5'b11011;
  /* fppowbf16.vhdl:736:28  */
  assign n6486 = x == 5'b11100;
  /* fppowbf16.vhdl:737:28  */
  assign n6489 = x == 5'b11101;
  /* fppowbf16.vhdl:738:28  */
  assign n6492 = x == 5'b11110;
  /* fppowbf16.vhdl:739:28  */
  assign n6495 = x == 5'b11111;
  assign n6497 = {n6495, n6492, n6489, n6486, n6483, n6480, n6477, n6474, n6471, n6468, n6465, n6462, n6459, n6456, n6453, n6450, n6447, n6444, n6441, n6438, n6435, n6432, n6429, n6426, n6423, n6420, n6417, n6414, n6411, n6408, n6405, n6402};
  /* fppowbf16.vhdl:707:4  */
  always @*
    case (n6497)
      32'b10000000000000000000000000000000: n6498 = 18'b101010111110011010;
      32'b01000000000000000000000000000000: n6498 = 18'b101001100101101100;
      32'b00100000000000000000000000000000: n6498 = 18'b101000001100111110;
      32'b00010000000000000000000000000000: n6498 = 18'b100110110100001111;
      32'b00001000000000000000000000000000: n6498 = 18'b100101011011100001;
      32'b00000100000000000000000000000000: n6498 = 18'b100100000010110011;
      32'b00000010000000000000000000000000: n6498 = 18'b100010101010000101;
      32'b00000001000000000000000000000000: n6498 = 18'b100001010001010110;
      32'b00000000100000000000000000000000: n6498 = 18'b011111111000101000;
      32'b00000000010000000000000000000000: n6498 = 18'b011110011111111010;
      32'b00000000001000000000000000000000: n6498 = 18'b011101000111001011;
      32'b00000000000100000000000000000000: n6498 = 18'b011011101110011101;
      32'b00000000000010000000000000000000: n6498 = 18'b011010010101101111;
      32'b00000000000001000000000000000000: n6498 = 18'b011000111101000001;
      32'b00000000000000100000000000000000: n6498 = 18'b010111100100010010;
      32'b00000000000000010000000000000000: n6498 = 18'b010110001011100100;
      32'b00000000000000001000000000000000: n6498 = 18'b010100110010110110;
      32'b00000000000000000100000000000000: n6498 = 18'b010011011010001000;
      32'b00000000000000000010000000000000: n6498 = 18'b010010000001011001;
      32'b00000000000000000001000000000000: n6498 = 18'b010000101000101011;
      32'b00000000000000000000100000000000: n6498 = 18'b001111001111111101;
      32'b00000000000000000000010000000000: n6498 = 18'b001101110111001111;
      32'b00000000000000000000001000000000: n6498 = 18'b001100011110100000;
      32'b00000000000000000000000100000000: n6498 = 18'b001011000101110010;
      32'b00000000000000000000000010000000: n6498 = 18'b001001101101000100;
      32'b00000000000000000000000001000000: n6498 = 18'b001000010100010110;
      32'b00000000000000000000000000100000: n6498 = 18'b000110111011100111;
      32'b00000000000000000000000000010000: n6498 = 18'b000101100010111001;
      32'b00000000000000000000000000001000: n6498 = 18'b000100001010001011;
      32'b00000000000000000000000000000100: n6498 = 18'b000010110001011101;
      32'b00000000000000000000000000000010: n6498 = 18'b000001011000101110;
      32'b00000000000000000000000000000001: n6498 = 18'b000000000000000000;
      default: n6498 = 18'bX;
    endcase
endmodule

module intadder_12_freq500_uid87
  (input  clk,
   input  [11:0] x,
   input  [11:0] y,
   input  cin,
   output [11:0] r);
  wire [11:0] rtmp;
  wire [11:0] x_d1;
  wire [11:0] y_d1;
  wire cin_d1;
  wire cin_d2;
  wire cin_d3;
  wire cin_d4;
  wire cin_d5;
  wire cin_d6;
  wire cin_d7;
  wire cin_d8;
  wire cin_d9;
  wire cin_d10;
  wire cin_d11;
  wire cin_d12;
  wire cin_d13;
  wire cin_d14;
  wire cin_d15;
  wire cin_d16;
  wire [11:0] n6378;
  wire [11:0] n6379;
  wire [11:0] n6380;
  reg [11:0] n6381;
  reg [11:0] n6382;
  reg n6383;
  reg n6384;
  reg n6385;
  reg n6386;
  reg n6387;
  reg n6388;
  reg n6389;
  reg n6390;
  reg n6391;
  reg n6392;
  reg n6393;
  reg n6394;
  reg n6395;
  reg n6396;
  reg n6397;
  reg n6398;
  assign r = rtmp; //(module output)
  /* fppowbf16.vhdl:4070:8  */
  assign rtmp = n6380; // (signal)
  /* fppowbf16.vhdl:4072:8  */
  assign x_d1 = n6381; // (signal)
  /* fppowbf16.vhdl:4074:8  */
  assign y_d1 = n6382; // (signal)
  /* fppowbf16.vhdl:4076:8  */
  assign cin_d1 = n6383; // (signal)
  /* fppowbf16.vhdl:4076:16  */
  assign cin_d2 = n6384; // (signal)
  /* fppowbf16.vhdl:4076:24  */
  assign cin_d3 = n6385; // (signal)
  /* fppowbf16.vhdl:4076:32  */
  assign cin_d4 = n6386; // (signal)
  /* fppowbf16.vhdl:4076:40  */
  assign cin_d5 = n6387; // (signal)
  /* fppowbf16.vhdl:4076:48  */
  assign cin_d6 = n6388; // (signal)
  /* fppowbf16.vhdl:4076:56  */
  assign cin_d7 = n6389; // (signal)
  /* fppowbf16.vhdl:4076:64  */
  assign cin_d8 = n6390; // (signal)
  /* fppowbf16.vhdl:4076:72  */
  assign cin_d9 = n6391; // (signal)
  /* fppowbf16.vhdl:4076:80  */
  assign cin_d10 = n6392; // (signal)
  /* fppowbf16.vhdl:4076:89  */
  assign cin_d11 = n6393; // (signal)
  /* fppowbf16.vhdl:4076:98  */
  assign cin_d12 = n6394; // (signal)
  /* fppowbf16.vhdl:4076:107  */
  assign cin_d13 = n6395; // (signal)
  /* fppowbf16.vhdl:4076:116  */
  assign cin_d14 = n6396; // (signal)
  /* fppowbf16.vhdl:4076:125  */
  assign cin_d15 = n6397; // (signal)
  /* fppowbf16.vhdl:4076:134  */
  assign cin_d16 = n6398; // (signal)
  /* fppowbf16.vhdl:4102:17  */
  assign n6378 = x_d1 + y_d1;
  /* fppowbf16.vhdl:4102:24  */
  assign n6379 = {11'b0, cin_d16};  //  uext
  /* fppowbf16.vhdl:4102:24  */
  assign n6380 = n6378 + n6379;
  /* fppowbf16.vhdl:4081:10  */
  always @(posedge clk)
    n6381 <= x;
  /* fppowbf16.vhdl:4081:10  */
  always @(posedge clk)
    n6382 <= y;
  /* fppowbf16.vhdl:4081:10  */
  always @(posedge clk)
    n6383 <= cin;
  /* fppowbf16.vhdl:4081:10  */
  always @(posedge clk)
    n6384 <= cin_d1;
  /* fppowbf16.vhdl:4081:10  */
  always @(posedge clk)
    n6385 <= cin_d2;
  /* fppowbf16.vhdl:4081:10  */
  always @(posedge clk)
    n6386 <= cin_d3;
  /* fppowbf16.vhdl:4081:10  */
  always @(posedge clk)
    n6387 <= cin_d4;
  /* fppowbf16.vhdl:4081:10  */
  always @(posedge clk)
    n6388 <= cin_d5;
  /* fppowbf16.vhdl:4081:10  */
  always @(posedge clk)
    n6389 <= cin_d6;
  /* fppowbf16.vhdl:4081:10  */
  always @(posedge clk)
    n6390 <= cin_d7;
  /* fppowbf16.vhdl:4081:10  */
  always @(posedge clk)
    n6391 <= cin_d8;
  /* fppowbf16.vhdl:4081:10  */
  always @(posedge clk)
    n6392 <= cin_d9;
  /* fppowbf16.vhdl:4081:10  */
  always @(posedge clk)
    n6393 <= cin_d10;
  /* fppowbf16.vhdl:4081:10  */
  always @(posedge clk)
    n6394 <= cin_d11;
  /* fppowbf16.vhdl:4081:10  */
  always @(posedge clk)
    n6395 <= cin_d12;
  /* fppowbf16.vhdl:4081:10  */
  always @(posedge clk)
    n6396 <= cin_d13;
  /* fppowbf16.vhdl:4081:10  */
  always @(posedge clk)
    n6397 <= cin_d14;
  /* fppowbf16.vhdl:4081:10  */
  always @(posedge clk)
    n6398 <= cin_d15;
endmodule

module fixrealkcm_freq500_uid77_t1_freq500_uid83
  (input  [4:0] x,
   output [6:0] y);
  wire [6:0] y0;
  wire [6:0] y1;
  wire n6258;
  wire n6261;
  wire n6264;
  wire n6267;
  wire n6270;
  wire n6273;
  wire n6276;
  wire n6279;
  wire n6282;
  wire n6285;
  wire n6288;
  wire n6291;
  wire n6294;
  wire n6297;
  wire n6300;
  wire n6303;
  wire n6306;
  wire n6309;
  wire n6312;
  wire n6315;
  wire n6318;
  wire n6321;
  wire n6324;
  wire n6327;
  wire n6330;
  wire n6333;
  wire n6336;
  wire n6339;
  wire n6342;
  wire n6345;
  wire n6348;
  wire n6351;
  wire [31:0] n6353;
  reg [6:0] n6354;
  assign y = y1; //(module output)
  /* fppowbf16.vhdl:630:8  */
  assign y0 = n6354; // (signal)
  /* fppowbf16.vhdl:632:8  */
  assign y1 = y0; // (signal)
  /* fppowbf16.vhdl:636:17  */
  assign n6258 = x == 5'b00000;
  /* fppowbf16.vhdl:637:17  */
  assign n6261 = x == 5'b00001;
  /* fppowbf16.vhdl:638:17  */
  assign n6264 = x == 5'b00010;
  /* fppowbf16.vhdl:639:17  */
  assign n6267 = x == 5'b00011;
  /* fppowbf16.vhdl:640:17  */
  assign n6270 = x == 5'b00100;
  /* fppowbf16.vhdl:641:17  */
  assign n6273 = x == 5'b00101;
  /* fppowbf16.vhdl:642:17  */
  assign n6276 = x == 5'b00110;
  /* fppowbf16.vhdl:643:17  */
  assign n6279 = x == 5'b00111;
  /* fppowbf16.vhdl:644:17  */
  assign n6282 = x == 5'b01000;
  /* fppowbf16.vhdl:645:17  */
  assign n6285 = x == 5'b01001;
  /* fppowbf16.vhdl:646:17  */
  assign n6288 = x == 5'b01010;
  /* fppowbf16.vhdl:647:17  */
  assign n6291 = x == 5'b01011;
  /* fppowbf16.vhdl:648:17  */
  assign n6294 = x == 5'b01100;
  /* fppowbf16.vhdl:649:17  */
  assign n6297 = x == 5'b01101;
  /* fppowbf16.vhdl:650:17  */
  assign n6300 = x == 5'b01110;
  /* fppowbf16.vhdl:651:17  */
  assign n6303 = x == 5'b01111;
  /* fppowbf16.vhdl:652:17  */
  assign n6306 = x == 5'b10000;
  /* fppowbf16.vhdl:653:17  */
  assign n6309 = x == 5'b10001;
  /* fppowbf16.vhdl:654:17  */
  assign n6312 = x == 5'b10010;
  /* fppowbf16.vhdl:655:17  */
  assign n6315 = x == 5'b10011;
  /* fppowbf16.vhdl:656:17  */
  assign n6318 = x == 5'b10100;
  /* fppowbf16.vhdl:657:17  */
  assign n6321 = x == 5'b10101;
  /* fppowbf16.vhdl:658:17  */
  assign n6324 = x == 5'b10110;
  /* fppowbf16.vhdl:659:17  */
  assign n6327 = x == 5'b10111;
  /* fppowbf16.vhdl:660:17  */
  assign n6330 = x == 5'b11000;
  /* fppowbf16.vhdl:661:17  */
  assign n6333 = x == 5'b11001;
  /* fppowbf16.vhdl:662:17  */
  assign n6336 = x == 5'b11010;
  /* fppowbf16.vhdl:663:17  */
  assign n6339 = x == 5'b11011;
  /* fppowbf16.vhdl:664:17  */
  assign n6342 = x == 5'b11100;
  /* fppowbf16.vhdl:665:17  */
  assign n6345 = x == 5'b11101;
  /* fppowbf16.vhdl:666:17  */
  assign n6348 = x == 5'b11110;
  /* fppowbf16.vhdl:667:17  */
  assign n6351 = x == 5'b11111;
  assign n6353 = {n6351, n6348, n6345, n6342, n6339, n6336, n6333, n6330, n6327, n6324, n6321, n6318, n6315, n6312, n6309, n6306, n6303, n6300, n6297, n6294, n6291, n6288, n6285, n6282, n6279, n6276, n6273, n6270, n6267, n6264, n6261, n6258};
  /* fppowbf16.vhdl:635:4  */
  always @*
    case (n6353)
      32'b10000000000000000000000000000000: n6354 = 7'b1011001;
      32'b01000000000000000000000000000000: n6354 = 7'b1010111;
      32'b00100000000000000000000000000000: n6354 = 7'b1010100;
      32'b00010000000000000000000000000000: n6354 = 7'b1010001;
      32'b00001000000000000000000000000000: n6354 = 7'b1001110;
      32'b00000100000000000000000000000000: n6354 = 7'b1001011;
      32'b00000010000000000000000000000000: n6354 = 7'b1001000;
      32'b00000001000000000000000000000000: n6354 = 7'b1000101;
      32'b00000000100000000000000000000000: n6354 = 7'b1000010;
      32'b00000000010000000000000000000000: n6354 = 7'b0111111;
      32'b00000000001000000000000000000000: n6354 = 7'b0111101;
      32'b00000000000100000000000000000000: n6354 = 7'b0111010;
      32'b00000000000010000000000000000000: n6354 = 7'b0110111;
      32'b00000000000001000000000000000000: n6354 = 7'b0110100;
      32'b00000000000000100000000000000000: n6354 = 7'b0110001;
      32'b00000000000000010000000000000000: n6354 = 7'b0101110;
      32'b00000000000000001000000000000000: n6354 = 7'b0101011;
      32'b00000000000000000100000000000000: n6354 = 7'b0101000;
      32'b00000000000000000010000000000000: n6354 = 7'b0100110;
      32'b00000000000000000001000000000000: n6354 = 7'b0100011;
      32'b00000000000000000000100000000000: n6354 = 7'b0100000;
      32'b00000000000000000000010000000000: n6354 = 7'b0011101;
      32'b00000000000000000000001000000000: n6354 = 7'b0011010;
      32'b00000000000000000000000100000000: n6354 = 7'b0010111;
      32'b00000000000000000000000010000000: n6354 = 7'b0010100;
      32'b00000000000000000000000001000000: n6354 = 7'b0010001;
      32'b00000000000000000000000000100000: n6354 = 7'b0001110;
      32'b00000000000000000000000000010000: n6354 = 7'b0001100;
      32'b00000000000000000000000000001000: n6354 = 7'b0001001;
      32'b00000000000000000000000000000100: n6354 = 7'b0000110;
      32'b00000000000000000000000000000010: n6354 = 7'b0000011;
      32'b00000000000000000000000000000001: n6354 = 7'b0000000;
      default: n6354 = 7'bX;
    endcase
endmodule

module fixrealkcm_freq500_uid77_t0_freq500_uid80
  (input  [4:0] x,
   output [11:0] y);
  wire [11:0] y0;
  wire [11:0] y1;
  wire n6158;
  wire n6161;
  wire n6164;
  wire n6167;
  wire n6170;
  wire n6173;
  wire n6176;
  wire n6179;
  wire n6182;
  wire n6185;
  wire n6188;
  wire n6191;
  wire n6194;
  wire n6197;
  wire n6200;
  wire n6203;
  wire n6206;
  wire n6209;
  wire n6212;
  wire n6215;
  wire n6218;
  wire n6221;
  wire n6224;
  wire n6227;
  wire n6230;
  wire n6233;
  wire n6236;
  wire n6239;
  wire n6242;
  wire n6245;
  wire n6248;
  wire n6251;
  wire [31:0] n6253;
  reg [11:0] n6254;
  assign y = y1; //(module output)
  /* fppowbf16.vhdl:558:8  */
  assign y0 = n6254; // (signal)
  /* fppowbf16.vhdl:560:8  */
  assign y1 = y0; // (signal)
  /* fppowbf16.vhdl:564:22  */
  assign n6158 = x == 5'b00000;
  /* fppowbf16.vhdl:565:22  */
  assign n6161 = x == 5'b00001;
  /* fppowbf16.vhdl:566:22  */
  assign n6164 = x == 5'b00010;
  /* fppowbf16.vhdl:567:22  */
  assign n6167 = x == 5'b00011;
  /* fppowbf16.vhdl:568:22  */
  assign n6170 = x == 5'b00100;
  /* fppowbf16.vhdl:569:22  */
  assign n6173 = x == 5'b00101;
  /* fppowbf16.vhdl:570:22  */
  assign n6176 = x == 5'b00110;
  /* fppowbf16.vhdl:571:22  */
  assign n6179 = x == 5'b00111;
  /* fppowbf16.vhdl:572:22  */
  assign n6182 = x == 5'b01000;
  /* fppowbf16.vhdl:573:22  */
  assign n6185 = x == 5'b01001;
  /* fppowbf16.vhdl:574:22  */
  assign n6188 = x == 5'b01010;
  /* fppowbf16.vhdl:575:22  */
  assign n6191 = x == 5'b01011;
  /* fppowbf16.vhdl:576:22  */
  assign n6194 = x == 5'b01100;
  /* fppowbf16.vhdl:577:22  */
  assign n6197 = x == 5'b01101;
  /* fppowbf16.vhdl:578:22  */
  assign n6200 = x == 5'b01110;
  /* fppowbf16.vhdl:579:22  */
  assign n6203 = x == 5'b01111;
  /* fppowbf16.vhdl:580:22  */
  assign n6206 = x == 5'b10000;
  /* fppowbf16.vhdl:581:22  */
  assign n6209 = x == 5'b10001;
  /* fppowbf16.vhdl:582:22  */
  assign n6212 = x == 5'b10010;
  /* fppowbf16.vhdl:583:22  */
  assign n6215 = x == 5'b10011;
  /* fppowbf16.vhdl:584:22  */
  assign n6218 = x == 5'b10100;
  /* fppowbf16.vhdl:585:22  */
  assign n6221 = x == 5'b10101;
  /* fppowbf16.vhdl:586:22  */
  assign n6224 = x == 5'b10110;
  /* fppowbf16.vhdl:587:22  */
  assign n6227 = x == 5'b10111;
  /* fppowbf16.vhdl:588:22  */
  assign n6230 = x == 5'b11000;
  /* fppowbf16.vhdl:589:22  */
  assign n6233 = x == 5'b11001;
  /* fppowbf16.vhdl:590:22  */
  assign n6236 = x == 5'b11010;
  /* fppowbf16.vhdl:591:22  */
  assign n6239 = x == 5'b11011;
  /* fppowbf16.vhdl:592:22  */
  assign n6242 = x == 5'b11100;
  /* fppowbf16.vhdl:593:22  */
  assign n6245 = x == 5'b11101;
  /* fppowbf16.vhdl:594:22  */
  assign n6248 = x == 5'b11110;
  /* fppowbf16.vhdl:595:22  */
  assign n6251 = x == 5'b11111;
  assign n6253 = {n6251, n6248, n6245, n6242, n6239, n6236, n6233, n6230, n6227, n6224, n6221, n6218, n6215, n6212, n6209, n6206, n6203, n6200, n6197, n6194, n6191, n6188, n6185, n6182, n6179, n6176, n6173, n6170, n6167, n6164, n6161, n6158};
  /* fppowbf16.vhdl:563:4  */
  always @*
    case (n6253)
      32'b10000000000000000000000000000000: n6254 = 12'b101100110110;
      32'b01000000000000000000000000000000: n6254 = 12'b101011011010;
      32'b00100000000000000000000000000000: n6254 = 12'b101001111110;
      32'b00010000000000000000000000000000: n6254 = 12'b101000100001;
      32'b00001000000000000000000000000000: n6254 = 12'b100111000101;
      32'b00000100000000000000000000000000: n6254 = 12'b100101101001;
      32'b00000010000000000000000000000000: n6254 = 12'b100100001100;
      32'b00000001000000000000000000000000: n6254 = 12'b100010110000;
      32'b00000000100000000000000000000000: n6254 = 12'b100001010100;
      32'b00000000010000000000000000000000: n6254 = 12'b011111110111;
      32'b00000000001000000000000000000000: n6254 = 12'b011110011011;
      32'b00000000000100000000000000000000: n6254 = 12'b011100111111;
      32'b00000000000010000000000000000000: n6254 = 12'b011011100010;
      32'b00000000000001000000000000000000: n6254 = 12'b011010000110;
      32'b00000000000000100000000000000000: n6254 = 12'b011000101010;
      32'b00000000000000010000000000000000: n6254 = 12'b010111001101;
      32'b00000000000000001000000000000000: n6254 = 12'b010101110001;
      32'b00000000000000000100000000000000: n6254 = 12'b010100010101;
      32'b00000000000000000010000000000000: n6254 = 12'b010010111000;
      32'b00000000000000000001000000000000: n6254 = 12'b010001011100;
      32'b00000000000000000000100000000000: n6254 = 12'b010000000000;
      32'b00000000000000000000010000000000: n6254 = 12'b001110100011;
      32'b00000000000000000000001000000000: n6254 = 12'b001101000111;
      32'b00000000000000000000000100000000: n6254 = 12'b001011101011;
      32'b00000000000000000000000010000000: n6254 = 12'b001010001110;
      32'b00000000000000000000000001000000: n6254 = 12'b001000110010;
      32'b00000000000000000000000000100000: n6254 = 12'b000111010110;
      32'b00000000000000000000000000010000: n6254 = 12'b000101111001;
      32'b00000000000000000000000000001000: n6254 = 12'b000100011101;
      32'b00000000000000000000000000000100: n6254 = 12'b000011000001;
      32'b00000000000000000000000000000010: n6254 = 12'b000001100100;
      32'b00000000000000000000000000000001: n6254 = 12'b000000001000;
      default: n6254 = 12'bX;
    endcase
endmodule

module fixfunctionbytable_freq500_uid104
  (input  [9:0] x,
   output [12:0] y);
  wire [12:0] y0;
  wire [12:0] y1;
  wire n3082;
  wire n3085;
  wire n3088;
  wire n3091;
  wire n3094;
  wire n3097;
  wire n3100;
  wire n3103;
  wire n3106;
  wire n3109;
  wire n3112;
  wire n3115;
  wire n3118;
  wire n3121;
  wire n3124;
  wire n3127;
  wire n3130;
  wire n3133;
  wire n3136;
  wire n3139;
  wire n3142;
  wire n3145;
  wire n3148;
  wire n3151;
  wire n3154;
  wire n3157;
  wire n3160;
  wire n3163;
  wire n3166;
  wire n3169;
  wire n3172;
  wire n3175;
  wire n3178;
  wire n3181;
  wire n3184;
  wire n3187;
  wire n3190;
  wire n3193;
  wire n3196;
  wire n3199;
  wire n3202;
  wire n3205;
  wire n3208;
  wire n3211;
  wire n3214;
  wire n3217;
  wire n3220;
  wire n3223;
  wire n3226;
  wire n3229;
  wire n3232;
  wire n3235;
  wire n3238;
  wire n3241;
  wire n3244;
  wire n3247;
  wire n3250;
  wire n3253;
  wire n3256;
  wire n3259;
  wire n3262;
  wire n3265;
  wire n3268;
  wire n3271;
  wire n3274;
  wire n3277;
  wire n3280;
  wire n3283;
  wire n3286;
  wire n3289;
  wire n3292;
  wire n3295;
  wire n3298;
  wire n3301;
  wire n3304;
  wire n3307;
  wire n3310;
  wire n3313;
  wire n3316;
  wire n3319;
  wire n3322;
  wire n3325;
  wire n3328;
  wire n3331;
  wire n3334;
  wire n3337;
  wire n3340;
  wire n3343;
  wire n3346;
  wire n3349;
  wire n3352;
  wire n3355;
  wire n3358;
  wire n3361;
  wire n3364;
  wire n3367;
  wire n3370;
  wire n3373;
  wire n3376;
  wire n3379;
  wire n3382;
  wire n3385;
  wire n3388;
  wire n3391;
  wire n3394;
  wire n3397;
  wire n3400;
  wire n3403;
  wire n3406;
  wire n3409;
  wire n3412;
  wire n3415;
  wire n3418;
  wire n3421;
  wire n3424;
  wire n3427;
  wire n3430;
  wire n3433;
  wire n3436;
  wire n3439;
  wire n3442;
  wire n3445;
  wire n3448;
  wire n3451;
  wire n3454;
  wire n3457;
  wire n3460;
  wire n3463;
  wire n3466;
  wire n3469;
  wire n3472;
  wire n3475;
  wire n3478;
  wire n3481;
  wire n3484;
  wire n3487;
  wire n3490;
  wire n3493;
  wire n3496;
  wire n3499;
  wire n3502;
  wire n3505;
  wire n3508;
  wire n3511;
  wire n3514;
  wire n3517;
  wire n3520;
  wire n3523;
  wire n3526;
  wire n3529;
  wire n3532;
  wire n3535;
  wire n3538;
  wire n3541;
  wire n3544;
  wire n3547;
  wire n3550;
  wire n3553;
  wire n3556;
  wire n3559;
  wire n3562;
  wire n3565;
  wire n3568;
  wire n3571;
  wire n3574;
  wire n3577;
  wire n3580;
  wire n3583;
  wire n3586;
  wire n3589;
  wire n3592;
  wire n3595;
  wire n3598;
  wire n3601;
  wire n3604;
  wire n3607;
  wire n3610;
  wire n3613;
  wire n3616;
  wire n3619;
  wire n3622;
  wire n3625;
  wire n3628;
  wire n3631;
  wire n3634;
  wire n3637;
  wire n3640;
  wire n3643;
  wire n3646;
  wire n3649;
  wire n3652;
  wire n3655;
  wire n3658;
  wire n3661;
  wire n3664;
  wire n3667;
  wire n3670;
  wire n3673;
  wire n3676;
  wire n3679;
  wire n3682;
  wire n3685;
  wire n3688;
  wire n3691;
  wire n3694;
  wire n3697;
  wire n3700;
  wire n3703;
  wire n3706;
  wire n3709;
  wire n3712;
  wire n3715;
  wire n3718;
  wire n3721;
  wire n3724;
  wire n3727;
  wire n3730;
  wire n3733;
  wire n3736;
  wire n3739;
  wire n3742;
  wire n3745;
  wire n3748;
  wire n3751;
  wire n3754;
  wire n3757;
  wire n3760;
  wire n3763;
  wire n3766;
  wire n3769;
  wire n3772;
  wire n3775;
  wire n3778;
  wire n3781;
  wire n3784;
  wire n3787;
  wire n3790;
  wire n3793;
  wire n3796;
  wire n3799;
  wire n3802;
  wire n3805;
  wire n3808;
  wire n3811;
  wire n3814;
  wire n3817;
  wire n3820;
  wire n3823;
  wire n3826;
  wire n3829;
  wire n3832;
  wire n3835;
  wire n3838;
  wire n3841;
  wire n3844;
  wire n3847;
  wire n3850;
  wire n3853;
  wire n3856;
  wire n3859;
  wire n3862;
  wire n3865;
  wire n3868;
  wire n3871;
  wire n3874;
  wire n3877;
  wire n3880;
  wire n3883;
  wire n3886;
  wire n3889;
  wire n3892;
  wire n3895;
  wire n3898;
  wire n3901;
  wire n3904;
  wire n3907;
  wire n3910;
  wire n3913;
  wire n3916;
  wire n3919;
  wire n3922;
  wire n3925;
  wire n3928;
  wire n3931;
  wire n3934;
  wire n3937;
  wire n3940;
  wire n3943;
  wire n3946;
  wire n3949;
  wire n3952;
  wire n3955;
  wire n3958;
  wire n3961;
  wire n3964;
  wire n3967;
  wire n3970;
  wire n3973;
  wire n3976;
  wire n3979;
  wire n3982;
  wire n3985;
  wire n3988;
  wire n3991;
  wire n3994;
  wire n3997;
  wire n4000;
  wire n4003;
  wire n4006;
  wire n4009;
  wire n4012;
  wire n4015;
  wire n4018;
  wire n4021;
  wire n4024;
  wire n4027;
  wire n4030;
  wire n4033;
  wire n4036;
  wire n4039;
  wire n4042;
  wire n4045;
  wire n4048;
  wire n4051;
  wire n4054;
  wire n4057;
  wire n4060;
  wire n4063;
  wire n4066;
  wire n4069;
  wire n4072;
  wire n4075;
  wire n4078;
  wire n4081;
  wire n4084;
  wire n4087;
  wire n4090;
  wire n4093;
  wire n4096;
  wire n4099;
  wire n4102;
  wire n4105;
  wire n4108;
  wire n4111;
  wire n4114;
  wire n4117;
  wire n4120;
  wire n4123;
  wire n4126;
  wire n4129;
  wire n4132;
  wire n4135;
  wire n4138;
  wire n4141;
  wire n4144;
  wire n4147;
  wire n4150;
  wire n4153;
  wire n4156;
  wire n4159;
  wire n4162;
  wire n4165;
  wire n4168;
  wire n4171;
  wire n4174;
  wire n4177;
  wire n4180;
  wire n4183;
  wire n4186;
  wire n4189;
  wire n4192;
  wire n4195;
  wire n4198;
  wire n4201;
  wire n4204;
  wire n4207;
  wire n4210;
  wire n4213;
  wire n4216;
  wire n4219;
  wire n4222;
  wire n4225;
  wire n4228;
  wire n4231;
  wire n4234;
  wire n4237;
  wire n4240;
  wire n4243;
  wire n4246;
  wire n4249;
  wire n4252;
  wire n4255;
  wire n4258;
  wire n4261;
  wire n4264;
  wire n4267;
  wire n4270;
  wire n4273;
  wire n4276;
  wire n4279;
  wire n4282;
  wire n4285;
  wire n4288;
  wire n4291;
  wire n4294;
  wire n4297;
  wire n4300;
  wire n4303;
  wire n4306;
  wire n4309;
  wire n4312;
  wire n4315;
  wire n4318;
  wire n4321;
  wire n4324;
  wire n4327;
  wire n4330;
  wire n4333;
  wire n4336;
  wire n4339;
  wire n4342;
  wire n4345;
  wire n4348;
  wire n4351;
  wire n4354;
  wire n4357;
  wire n4360;
  wire n4363;
  wire n4366;
  wire n4369;
  wire n4372;
  wire n4375;
  wire n4378;
  wire n4381;
  wire n4384;
  wire n4387;
  wire n4390;
  wire n4393;
  wire n4396;
  wire n4399;
  wire n4402;
  wire n4405;
  wire n4408;
  wire n4411;
  wire n4414;
  wire n4417;
  wire n4420;
  wire n4423;
  wire n4426;
  wire n4429;
  wire n4432;
  wire n4435;
  wire n4438;
  wire n4441;
  wire n4444;
  wire n4447;
  wire n4450;
  wire n4453;
  wire n4456;
  wire n4459;
  wire n4462;
  wire n4465;
  wire n4468;
  wire n4471;
  wire n4474;
  wire n4477;
  wire n4480;
  wire n4483;
  wire n4486;
  wire n4489;
  wire n4492;
  wire n4495;
  wire n4498;
  wire n4501;
  wire n4504;
  wire n4507;
  wire n4510;
  wire n4513;
  wire n4516;
  wire n4519;
  wire n4522;
  wire n4525;
  wire n4528;
  wire n4531;
  wire n4534;
  wire n4537;
  wire n4540;
  wire n4543;
  wire n4546;
  wire n4549;
  wire n4552;
  wire n4555;
  wire n4558;
  wire n4561;
  wire n4564;
  wire n4567;
  wire n4570;
  wire n4573;
  wire n4576;
  wire n4579;
  wire n4582;
  wire n4585;
  wire n4588;
  wire n4591;
  wire n4594;
  wire n4597;
  wire n4600;
  wire n4603;
  wire n4606;
  wire n4609;
  wire n4612;
  wire n4615;
  wire n4618;
  wire n4621;
  wire n4624;
  wire n4627;
  wire n4630;
  wire n4633;
  wire n4636;
  wire n4639;
  wire n4642;
  wire n4645;
  wire n4648;
  wire n4651;
  wire n4654;
  wire n4657;
  wire n4660;
  wire n4663;
  wire n4666;
  wire n4669;
  wire n4672;
  wire n4675;
  wire n4678;
  wire n4681;
  wire n4684;
  wire n4687;
  wire n4690;
  wire n4693;
  wire n4696;
  wire n4699;
  wire n4702;
  wire n4705;
  wire n4708;
  wire n4711;
  wire n4714;
  wire n4717;
  wire n4720;
  wire n4723;
  wire n4726;
  wire n4729;
  wire n4732;
  wire n4735;
  wire n4738;
  wire n4741;
  wire n4744;
  wire n4747;
  wire n4750;
  wire n4753;
  wire n4756;
  wire n4759;
  wire n4762;
  wire n4765;
  wire n4768;
  wire n4771;
  wire n4774;
  wire n4777;
  wire n4780;
  wire n4783;
  wire n4786;
  wire n4789;
  wire n4792;
  wire n4795;
  wire n4798;
  wire n4801;
  wire n4804;
  wire n4807;
  wire n4810;
  wire n4813;
  wire n4816;
  wire n4819;
  wire n4822;
  wire n4825;
  wire n4828;
  wire n4831;
  wire n4834;
  wire n4837;
  wire n4840;
  wire n4843;
  wire n4846;
  wire n4849;
  wire n4852;
  wire n4855;
  wire n4858;
  wire n4861;
  wire n4864;
  wire n4867;
  wire n4870;
  wire n4873;
  wire n4876;
  wire n4879;
  wire n4882;
  wire n4885;
  wire n4888;
  wire n4891;
  wire n4894;
  wire n4897;
  wire n4900;
  wire n4903;
  wire n4906;
  wire n4909;
  wire n4912;
  wire n4915;
  wire n4918;
  wire n4921;
  wire n4924;
  wire n4927;
  wire n4930;
  wire n4933;
  wire n4936;
  wire n4939;
  wire n4942;
  wire n4945;
  wire n4948;
  wire n4951;
  wire n4954;
  wire n4957;
  wire n4960;
  wire n4963;
  wire n4966;
  wire n4969;
  wire n4972;
  wire n4975;
  wire n4978;
  wire n4981;
  wire n4984;
  wire n4987;
  wire n4990;
  wire n4993;
  wire n4996;
  wire n4999;
  wire n5002;
  wire n5005;
  wire n5008;
  wire n5011;
  wire n5014;
  wire n5017;
  wire n5020;
  wire n5023;
  wire n5026;
  wire n5029;
  wire n5032;
  wire n5035;
  wire n5038;
  wire n5041;
  wire n5044;
  wire n5047;
  wire n5050;
  wire n5053;
  wire n5056;
  wire n5059;
  wire n5062;
  wire n5065;
  wire n5068;
  wire n5071;
  wire n5074;
  wire n5077;
  wire n5080;
  wire n5083;
  wire n5086;
  wire n5089;
  wire n5092;
  wire n5095;
  wire n5098;
  wire n5101;
  wire n5104;
  wire n5107;
  wire n5110;
  wire n5113;
  wire n5116;
  wire n5119;
  wire n5122;
  wire n5125;
  wire n5128;
  wire n5131;
  wire n5134;
  wire n5137;
  wire n5140;
  wire n5143;
  wire n5146;
  wire n5149;
  wire n5152;
  wire n5155;
  wire n5158;
  wire n5161;
  wire n5164;
  wire n5167;
  wire n5170;
  wire n5173;
  wire n5176;
  wire n5179;
  wire n5182;
  wire n5185;
  wire n5188;
  wire n5191;
  wire n5194;
  wire n5197;
  wire n5200;
  wire n5203;
  wire n5206;
  wire n5209;
  wire n5212;
  wire n5215;
  wire n5218;
  wire n5221;
  wire n5224;
  wire n5227;
  wire n5230;
  wire n5233;
  wire n5236;
  wire n5239;
  wire n5242;
  wire n5245;
  wire n5248;
  wire n5251;
  wire n5254;
  wire n5257;
  wire n5260;
  wire n5263;
  wire n5266;
  wire n5269;
  wire n5272;
  wire n5275;
  wire n5278;
  wire n5281;
  wire n5284;
  wire n5287;
  wire n5290;
  wire n5293;
  wire n5296;
  wire n5299;
  wire n5302;
  wire n5305;
  wire n5308;
  wire n5311;
  wire n5314;
  wire n5317;
  wire n5320;
  wire n5323;
  wire n5326;
  wire n5329;
  wire n5332;
  wire n5335;
  wire n5338;
  wire n5341;
  wire n5344;
  wire n5347;
  wire n5350;
  wire n5353;
  wire n5356;
  wire n5359;
  wire n5362;
  wire n5365;
  wire n5368;
  wire n5371;
  wire n5374;
  wire n5377;
  wire n5380;
  wire n5383;
  wire n5386;
  wire n5389;
  wire n5392;
  wire n5395;
  wire n5398;
  wire n5401;
  wire n5404;
  wire n5407;
  wire n5410;
  wire n5413;
  wire n5416;
  wire n5419;
  wire n5422;
  wire n5425;
  wire n5428;
  wire n5431;
  wire n5434;
  wire n5437;
  wire n5440;
  wire n5443;
  wire n5446;
  wire n5449;
  wire n5452;
  wire n5455;
  wire n5458;
  wire n5461;
  wire n5464;
  wire n5467;
  wire n5470;
  wire n5473;
  wire n5476;
  wire n5479;
  wire n5482;
  wire n5485;
  wire n5488;
  wire n5491;
  wire n5494;
  wire n5497;
  wire n5500;
  wire n5503;
  wire n5506;
  wire n5509;
  wire n5512;
  wire n5515;
  wire n5518;
  wire n5521;
  wire n5524;
  wire n5527;
  wire n5530;
  wire n5533;
  wire n5536;
  wire n5539;
  wire n5542;
  wire n5545;
  wire n5548;
  wire n5551;
  wire n5554;
  wire n5557;
  wire n5560;
  wire n5563;
  wire n5566;
  wire n5569;
  wire n5572;
  wire n5575;
  wire n5578;
  wire n5581;
  wire n5584;
  wire n5587;
  wire n5590;
  wire n5593;
  wire n5596;
  wire n5599;
  wire n5602;
  wire n5605;
  wire n5608;
  wire n5611;
  wire n5614;
  wire n5617;
  wire n5620;
  wire n5623;
  wire n5626;
  wire n5629;
  wire n5632;
  wire n5635;
  wire n5638;
  wire n5641;
  wire n5644;
  wire n5647;
  wire n5650;
  wire n5653;
  wire n5656;
  wire n5659;
  wire n5662;
  wire n5665;
  wire n5668;
  wire n5671;
  wire n5674;
  wire n5677;
  wire n5680;
  wire n5683;
  wire n5686;
  wire n5689;
  wire n5692;
  wire n5695;
  wire n5698;
  wire n5701;
  wire n5704;
  wire n5707;
  wire n5710;
  wire n5713;
  wire n5716;
  wire n5719;
  wire n5722;
  wire n5725;
  wire n5728;
  wire n5731;
  wire n5734;
  wire n5737;
  wire n5740;
  wire n5743;
  wire n5746;
  wire n5749;
  wire n5752;
  wire n5755;
  wire n5758;
  wire n5761;
  wire n5764;
  wire n5767;
  wire n5770;
  wire n5773;
  wire n5776;
  wire n5779;
  wire n5782;
  wire n5785;
  wire n5788;
  wire n5791;
  wire n5794;
  wire n5797;
  wire n5800;
  wire n5803;
  wire n5806;
  wire n5809;
  wire n5812;
  wire n5815;
  wire n5818;
  wire n5821;
  wire n5824;
  wire n5827;
  wire n5830;
  wire n5833;
  wire n5836;
  wire n5839;
  wire n5842;
  wire n5845;
  wire n5848;
  wire n5851;
  wire n5854;
  wire n5857;
  wire n5860;
  wire n5863;
  wire n5866;
  wire n5869;
  wire n5872;
  wire n5875;
  wire n5878;
  wire n5881;
  wire n5884;
  wire n5887;
  wire n5890;
  wire n5893;
  wire n5896;
  wire n5899;
  wire n5902;
  wire n5905;
  wire n5908;
  wire n5911;
  wire n5914;
  wire n5917;
  wire n5920;
  wire n5923;
  wire n5926;
  wire n5929;
  wire n5932;
  wire n5935;
  wire n5938;
  wire n5941;
  wire n5944;
  wire n5947;
  wire n5950;
  wire n5953;
  wire n5956;
  wire n5959;
  wire n5962;
  wire n5965;
  wire n5968;
  wire n5971;
  wire n5974;
  wire n5977;
  wire n5980;
  wire n5983;
  wire n5986;
  wire n5989;
  wire n5992;
  wire n5995;
  wire n5998;
  wire n6001;
  wire n6004;
  wire n6007;
  wire n6010;
  wire n6013;
  wire n6016;
  wire n6019;
  wire n6022;
  wire n6025;
  wire n6028;
  wire n6031;
  wire n6034;
  wire n6037;
  wire n6040;
  wire n6043;
  wire n6046;
  wire n6049;
  wire n6052;
  wire n6055;
  wire n6058;
  wire n6061;
  wire n6064;
  wire n6067;
  wire n6070;
  wire n6073;
  wire n6076;
  wire n6079;
  wire n6082;
  wire n6085;
  wire n6088;
  wire n6091;
  wire n6094;
  wire n6097;
  wire n6100;
  wire n6103;
  wire n6106;
  wire n6109;
  wire n6112;
  wire n6115;
  wire n6118;
  wire n6121;
  wire n6124;
  wire n6127;
  wire n6130;
  wire n6133;
  wire n6136;
  wire n6139;
  wire n6142;
  wire n6145;
  wire n6148;
  wire n6151;
  wire [1023:0] n6153;
  reg [12:0] n6154;
  assign y = y1; //(module output)
  /* fppowbf16.vhdl:824:8  */
  assign y0 = n6154; // (signal)
  /* fppowbf16.vhdl:826:8  */
  assign y1 = y0; // (signal)
  /* fppowbf16.vhdl:830:23  */
  assign n3082 = x == 10'b0000000000;
  /* fppowbf16.vhdl:831:23  */
  assign n3085 = x == 10'b0000000001;
  /* fppowbf16.vhdl:832:23  */
  assign n3088 = x == 10'b0000000010;
  /* fppowbf16.vhdl:833:23  */
  assign n3091 = x == 10'b0000000011;
  /* fppowbf16.vhdl:834:23  */
  assign n3094 = x == 10'b0000000100;
  /* fppowbf16.vhdl:835:23  */
  assign n3097 = x == 10'b0000000101;
  /* fppowbf16.vhdl:836:23  */
  assign n3100 = x == 10'b0000000110;
  /* fppowbf16.vhdl:837:23  */
  assign n3103 = x == 10'b0000000111;
  /* fppowbf16.vhdl:838:23  */
  assign n3106 = x == 10'b0000001000;
  /* fppowbf16.vhdl:839:23  */
  assign n3109 = x == 10'b0000001001;
  /* fppowbf16.vhdl:840:23  */
  assign n3112 = x == 10'b0000001010;
  /* fppowbf16.vhdl:841:23  */
  assign n3115 = x == 10'b0000001011;
  /* fppowbf16.vhdl:842:23  */
  assign n3118 = x == 10'b0000001100;
  /* fppowbf16.vhdl:843:23  */
  assign n3121 = x == 10'b0000001101;
  /* fppowbf16.vhdl:844:23  */
  assign n3124 = x == 10'b0000001110;
  /* fppowbf16.vhdl:845:23  */
  assign n3127 = x == 10'b0000001111;
  /* fppowbf16.vhdl:846:23  */
  assign n3130 = x == 10'b0000010000;
  /* fppowbf16.vhdl:847:23  */
  assign n3133 = x == 10'b0000010001;
  /* fppowbf16.vhdl:848:23  */
  assign n3136 = x == 10'b0000010010;
  /* fppowbf16.vhdl:849:23  */
  assign n3139 = x == 10'b0000010011;
  /* fppowbf16.vhdl:850:23  */
  assign n3142 = x == 10'b0000010100;
  /* fppowbf16.vhdl:851:23  */
  assign n3145 = x == 10'b0000010101;
  /* fppowbf16.vhdl:852:23  */
  assign n3148 = x == 10'b0000010110;
  /* fppowbf16.vhdl:853:23  */
  assign n3151 = x == 10'b0000010111;
  /* fppowbf16.vhdl:854:23  */
  assign n3154 = x == 10'b0000011000;
  /* fppowbf16.vhdl:855:23  */
  assign n3157 = x == 10'b0000011001;
  /* fppowbf16.vhdl:856:23  */
  assign n3160 = x == 10'b0000011010;
  /* fppowbf16.vhdl:857:23  */
  assign n3163 = x == 10'b0000011011;
  /* fppowbf16.vhdl:858:23  */
  assign n3166 = x == 10'b0000011100;
  /* fppowbf16.vhdl:859:23  */
  assign n3169 = x == 10'b0000011101;
  /* fppowbf16.vhdl:860:23  */
  assign n3172 = x == 10'b0000011110;
  /* fppowbf16.vhdl:861:23  */
  assign n3175 = x == 10'b0000011111;
  /* fppowbf16.vhdl:862:23  */
  assign n3178 = x == 10'b0000100000;
  /* fppowbf16.vhdl:863:23  */
  assign n3181 = x == 10'b0000100001;
  /* fppowbf16.vhdl:864:23  */
  assign n3184 = x == 10'b0000100010;
  /* fppowbf16.vhdl:865:23  */
  assign n3187 = x == 10'b0000100011;
  /* fppowbf16.vhdl:866:23  */
  assign n3190 = x == 10'b0000100100;
  /* fppowbf16.vhdl:867:23  */
  assign n3193 = x == 10'b0000100101;
  /* fppowbf16.vhdl:868:23  */
  assign n3196 = x == 10'b0000100110;
  /* fppowbf16.vhdl:869:23  */
  assign n3199 = x == 10'b0000100111;
  /* fppowbf16.vhdl:870:23  */
  assign n3202 = x == 10'b0000101000;
  /* fppowbf16.vhdl:871:23  */
  assign n3205 = x == 10'b0000101001;
  /* fppowbf16.vhdl:872:23  */
  assign n3208 = x == 10'b0000101010;
  /* fppowbf16.vhdl:873:23  */
  assign n3211 = x == 10'b0000101011;
  /* fppowbf16.vhdl:874:23  */
  assign n3214 = x == 10'b0000101100;
  /* fppowbf16.vhdl:875:23  */
  assign n3217 = x == 10'b0000101101;
  /* fppowbf16.vhdl:876:23  */
  assign n3220 = x == 10'b0000101110;
  /* fppowbf16.vhdl:877:23  */
  assign n3223 = x == 10'b0000101111;
  /* fppowbf16.vhdl:878:23  */
  assign n3226 = x == 10'b0000110000;
  /* fppowbf16.vhdl:879:23  */
  assign n3229 = x == 10'b0000110001;
  /* fppowbf16.vhdl:880:23  */
  assign n3232 = x == 10'b0000110010;
  /* fppowbf16.vhdl:881:23  */
  assign n3235 = x == 10'b0000110011;
  /* fppowbf16.vhdl:882:23  */
  assign n3238 = x == 10'b0000110100;
  /* fppowbf16.vhdl:883:23  */
  assign n3241 = x == 10'b0000110101;
  /* fppowbf16.vhdl:884:23  */
  assign n3244 = x == 10'b0000110110;
  /* fppowbf16.vhdl:885:23  */
  assign n3247 = x == 10'b0000110111;
  /* fppowbf16.vhdl:886:23  */
  assign n3250 = x == 10'b0000111000;
  /* fppowbf16.vhdl:887:23  */
  assign n3253 = x == 10'b0000111001;
  /* fppowbf16.vhdl:888:23  */
  assign n3256 = x == 10'b0000111010;
  /* fppowbf16.vhdl:889:23  */
  assign n3259 = x == 10'b0000111011;
  /* fppowbf16.vhdl:890:23  */
  assign n3262 = x == 10'b0000111100;
  /* fppowbf16.vhdl:891:23  */
  assign n3265 = x == 10'b0000111101;
  /* fppowbf16.vhdl:892:23  */
  assign n3268 = x == 10'b0000111110;
  /* fppowbf16.vhdl:893:23  */
  assign n3271 = x == 10'b0000111111;
  /* fppowbf16.vhdl:894:23  */
  assign n3274 = x == 10'b0001000000;
  /* fppowbf16.vhdl:895:23  */
  assign n3277 = x == 10'b0001000001;
  /* fppowbf16.vhdl:896:23  */
  assign n3280 = x == 10'b0001000010;
  /* fppowbf16.vhdl:897:23  */
  assign n3283 = x == 10'b0001000011;
  /* fppowbf16.vhdl:898:23  */
  assign n3286 = x == 10'b0001000100;
  /* fppowbf16.vhdl:899:23  */
  assign n3289 = x == 10'b0001000101;
  /* fppowbf16.vhdl:900:23  */
  assign n3292 = x == 10'b0001000110;
  /* fppowbf16.vhdl:901:23  */
  assign n3295 = x == 10'b0001000111;
  /* fppowbf16.vhdl:902:23  */
  assign n3298 = x == 10'b0001001000;
  /* fppowbf16.vhdl:903:23  */
  assign n3301 = x == 10'b0001001001;
  /* fppowbf16.vhdl:904:23  */
  assign n3304 = x == 10'b0001001010;
  /* fppowbf16.vhdl:905:23  */
  assign n3307 = x == 10'b0001001011;
  /* fppowbf16.vhdl:906:23  */
  assign n3310 = x == 10'b0001001100;
  /* fppowbf16.vhdl:907:23  */
  assign n3313 = x == 10'b0001001101;
  /* fppowbf16.vhdl:908:23  */
  assign n3316 = x == 10'b0001001110;
  /* fppowbf16.vhdl:909:23  */
  assign n3319 = x == 10'b0001001111;
  /* fppowbf16.vhdl:910:23  */
  assign n3322 = x == 10'b0001010000;
  /* fppowbf16.vhdl:911:23  */
  assign n3325 = x == 10'b0001010001;
  /* fppowbf16.vhdl:912:23  */
  assign n3328 = x == 10'b0001010010;
  /* fppowbf16.vhdl:913:23  */
  assign n3331 = x == 10'b0001010011;
  /* fppowbf16.vhdl:914:23  */
  assign n3334 = x == 10'b0001010100;
  /* fppowbf16.vhdl:915:23  */
  assign n3337 = x == 10'b0001010101;
  /* fppowbf16.vhdl:916:23  */
  assign n3340 = x == 10'b0001010110;
  /* fppowbf16.vhdl:917:23  */
  assign n3343 = x == 10'b0001010111;
  /* fppowbf16.vhdl:918:23  */
  assign n3346 = x == 10'b0001011000;
  /* fppowbf16.vhdl:919:23  */
  assign n3349 = x == 10'b0001011001;
  /* fppowbf16.vhdl:920:23  */
  assign n3352 = x == 10'b0001011010;
  /* fppowbf16.vhdl:921:23  */
  assign n3355 = x == 10'b0001011011;
  /* fppowbf16.vhdl:922:23  */
  assign n3358 = x == 10'b0001011100;
  /* fppowbf16.vhdl:923:23  */
  assign n3361 = x == 10'b0001011101;
  /* fppowbf16.vhdl:924:23  */
  assign n3364 = x == 10'b0001011110;
  /* fppowbf16.vhdl:925:23  */
  assign n3367 = x == 10'b0001011111;
  /* fppowbf16.vhdl:926:23  */
  assign n3370 = x == 10'b0001100000;
  /* fppowbf16.vhdl:927:23  */
  assign n3373 = x == 10'b0001100001;
  /* fppowbf16.vhdl:928:23  */
  assign n3376 = x == 10'b0001100010;
  /* fppowbf16.vhdl:929:23  */
  assign n3379 = x == 10'b0001100011;
  /* fppowbf16.vhdl:930:23  */
  assign n3382 = x == 10'b0001100100;
  /* fppowbf16.vhdl:931:23  */
  assign n3385 = x == 10'b0001100101;
  /* fppowbf16.vhdl:932:23  */
  assign n3388 = x == 10'b0001100110;
  /* fppowbf16.vhdl:933:23  */
  assign n3391 = x == 10'b0001100111;
  /* fppowbf16.vhdl:934:23  */
  assign n3394 = x == 10'b0001101000;
  /* fppowbf16.vhdl:935:23  */
  assign n3397 = x == 10'b0001101001;
  /* fppowbf16.vhdl:936:23  */
  assign n3400 = x == 10'b0001101010;
  /* fppowbf16.vhdl:937:23  */
  assign n3403 = x == 10'b0001101011;
  /* fppowbf16.vhdl:938:23  */
  assign n3406 = x == 10'b0001101100;
  /* fppowbf16.vhdl:939:23  */
  assign n3409 = x == 10'b0001101101;
  /* fppowbf16.vhdl:940:23  */
  assign n3412 = x == 10'b0001101110;
  /* fppowbf16.vhdl:941:23  */
  assign n3415 = x == 10'b0001101111;
  /* fppowbf16.vhdl:942:23  */
  assign n3418 = x == 10'b0001110000;
  /* fppowbf16.vhdl:943:23  */
  assign n3421 = x == 10'b0001110001;
  /* fppowbf16.vhdl:944:23  */
  assign n3424 = x == 10'b0001110010;
  /* fppowbf16.vhdl:945:23  */
  assign n3427 = x == 10'b0001110011;
  /* fppowbf16.vhdl:946:23  */
  assign n3430 = x == 10'b0001110100;
  /* fppowbf16.vhdl:947:23  */
  assign n3433 = x == 10'b0001110101;
  /* fppowbf16.vhdl:948:23  */
  assign n3436 = x == 10'b0001110110;
  /* fppowbf16.vhdl:949:23  */
  assign n3439 = x == 10'b0001110111;
  /* fppowbf16.vhdl:950:23  */
  assign n3442 = x == 10'b0001111000;
  /* fppowbf16.vhdl:951:23  */
  assign n3445 = x == 10'b0001111001;
  /* fppowbf16.vhdl:952:23  */
  assign n3448 = x == 10'b0001111010;
  /* fppowbf16.vhdl:953:23  */
  assign n3451 = x == 10'b0001111011;
  /* fppowbf16.vhdl:954:23  */
  assign n3454 = x == 10'b0001111100;
  /* fppowbf16.vhdl:955:23  */
  assign n3457 = x == 10'b0001111101;
  /* fppowbf16.vhdl:956:23  */
  assign n3460 = x == 10'b0001111110;
  /* fppowbf16.vhdl:957:23  */
  assign n3463 = x == 10'b0001111111;
  /* fppowbf16.vhdl:958:23  */
  assign n3466 = x == 10'b0010000000;
  /* fppowbf16.vhdl:959:23  */
  assign n3469 = x == 10'b0010000001;
  /* fppowbf16.vhdl:960:23  */
  assign n3472 = x == 10'b0010000010;
  /* fppowbf16.vhdl:961:23  */
  assign n3475 = x == 10'b0010000011;
  /* fppowbf16.vhdl:962:23  */
  assign n3478 = x == 10'b0010000100;
  /* fppowbf16.vhdl:963:23  */
  assign n3481 = x == 10'b0010000101;
  /* fppowbf16.vhdl:964:23  */
  assign n3484 = x == 10'b0010000110;
  /* fppowbf16.vhdl:965:23  */
  assign n3487 = x == 10'b0010000111;
  /* fppowbf16.vhdl:966:23  */
  assign n3490 = x == 10'b0010001000;
  /* fppowbf16.vhdl:967:23  */
  assign n3493 = x == 10'b0010001001;
  /* fppowbf16.vhdl:968:23  */
  assign n3496 = x == 10'b0010001010;
  /* fppowbf16.vhdl:969:23  */
  assign n3499 = x == 10'b0010001011;
  /* fppowbf16.vhdl:970:23  */
  assign n3502 = x == 10'b0010001100;
  /* fppowbf16.vhdl:971:23  */
  assign n3505 = x == 10'b0010001101;
  /* fppowbf16.vhdl:972:23  */
  assign n3508 = x == 10'b0010001110;
  /* fppowbf16.vhdl:973:23  */
  assign n3511 = x == 10'b0010001111;
  /* fppowbf16.vhdl:974:23  */
  assign n3514 = x == 10'b0010010000;
  /* fppowbf16.vhdl:975:23  */
  assign n3517 = x == 10'b0010010001;
  /* fppowbf16.vhdl:976:23  */
  assign n3520 = x == 10'b0010010010;
  /* fppowbf16.vhdl:977:23  */
  assign n3523 = x == 10'b0010010011;
  /* fppowbf16.vhdl:978:23  */
  assign n3526 = x == 10'b0010010100;
  /* fppowbf16.vhdl:979:23  */
  assign n3529 = x == 10'b0010010101;
  /* fppowbf16.vhdl:980:23  */
  assign n3532 = x == 10'b0010010110;
  /* fppowbf16.vhdl:981:23  */
  assign n3535 = x == 10'b0010010111;
  /* fppowbf16.vhdl:982:23  */
  assign n3538 = x == 10'b0010011000;
  /* fppowbf16.vhdl:983:23  */
  assign n3541 = x == 10'b0010011001;
  /* fppowbf16.vhdl:984:23  */
  assign n3544 = x == 10'b0010011010;
  /* fppowbf16.vhdl:985:23  */
  assign n3547 = x == 10'b0010011011;
  /* fppowbf16.vhdl:986:23  */
  assign n3550 = x == 10'b0010011100;
  /* fppowbf16.vhdl:987:23  */
  assign n3553 = x == 10'b0010011101;
  /* fppowbf16.vhdl:988:23  */
  assign n3556 = x == 10'b0010011110;
  /* fppowbf16.vhdl:989:23  */
  assign n3559 = x == 10'b0010011111;
  /* fppowbf16.vhdl:990:23  */
  assign n3562 = x == 10'b0010100000;
  /* fppowbf16.vhdl:991:23  */
  assign n3565 = x == 10'b0010100001;
  /* fppowbf16.vhdl:992:23  */
  assign n3568 = x == 10'b0010100010;
  /* fppowbf16.vhdl:993:23  */
  assign n3571 = x == 10'b0010100011;
  /* fppowbf16.vhdl:994:23  */
  assign n3574 = x == 10'b0010100100;
  /* fppowbf16.vhdl:995:23  */
  assign n3577 = x == 10'b0010100101;
  /* fppowbf16.vhdl:996:23  */
  assign n3580 = x == 10'b0010100110;
  /* fppowbf16.vhdl:997:23  */
  assign n3583 = x == 10'b0010100111;
  /* fppowbf16.vhdl:998:23  */
  assign n3586 = x == 10'b0010101000;
  /* fppowbf16.vhdl:999:23  */
  assign n3589 = x == 10'b0010101001;
  /* fppowbf16.vhdl:1000:23  */
  assign n3592 = x == 10'b0010101010;
  /* fppowbf16.vhdl:1001:23  */
  assign n3595 = x == 10'b0010101011;
  /* fppowbf16.vhdl:1002:23  */
  assign n3598 = x == 10'b0010101100;
  /* fppowbf16.vhdl:1003:23  */
  assign n3601 = x == 10'b0010101101;
  /* fppowbf16.vhdl:1004:23  */
  assign n3604 = x == 10'b0010101110;
  /* fppowbf16.vhdl:1005:23  */
  assign n3607 = x == 10'b0010101111;
  /* fppowbf16.vhdl:1006:23  */
  assign n3610 = x == 10'b0010110000;
  /* fppowbf16.vhdl:1007:23  */
  assign n3613 = x == 10'b0010110001;
  /* fppowbf16.vhdl:1008:23  */
  assign n3616 = x == 10'b0010110010;
  /* fppowbf16.vhdl:1009:23  */
  assign n3619 = x == 10'b0010110011;
  /* fppowbf16.vhdl:1010:23  */
  assign n3622 = x == 10'b0010110100;
  /* fppowbf16.vhdl:1011:23  */
  assign n3625 = x == 10'b0010110101;
  /* fppowbf16.vhdl:1012:23  */
  assign n3628 = x == 10'b0010110110;
  /* fppowbf16.vhdl:1013:23  */
  assign n3631 = x == 10'b0010110111;
  /* fppowbf16.vhdl:1014:23  */
  assign n3634 = x == 10'b0010111000;
  /* fppowbf16.vhdl:1015:23  */
  assign n3637 = x == 10'b0010111001;
  /* fppowbf16.vhdl:1016:23  */
  assign n3640 = x == 10'b0010111010;
  /* fppowbf16.vhdl:1017:23  */
  assign n3643 = x == 10'b0010111011;
  /* fppowbf16.vhdl:1018:23  */
  assign n3646 = x == 10'b0010111100;
  /* fppowbf16.vhdl:1019:23  */
  assign n3649 = x == 10'b0010111101;
  /* fppowbf16.vhdl:1020:23  */
  assign n3652 = x == 10'b0010111110;
  /* fppowbf16.vhdl:1021:23  */
  assign n3655 = x == 10'b0010111111;
  /* fppowbf16.vhdl:1022:23  */
  assign n3658 = x == 10'b0011000000;
  /* fppowbf16.vhdl:1023:23  */
  assign n3661 = x == 10'b0011000001;
  /* fppowbf16.vhdl:1024:23  */
  assign n3664 = x == 10'b0011000010;
  /* fppowbf16.vhdl:1025:23  */
  assign n3667 = x == 10'b0011000011;
  /* fppowbf16.vhdl:1026:23  */
  assign n3670 = x == 10'b0011000100;
  /* fppowbf16.vhdl:1027:23  */
  assign n3673 = x == 10'b0011000101;
  /* fppowbf16.vhdl:1028:23  */
  assign n3676 = x == 10'b0011000110;
  /* fppowbf16.vhdl:1029:23  */
  assign n3679 = x == 10'b0011000111;
  /* fppowbf16.vhdl:1030:23  */
  assign n3682 = x == 10'b0011001000;
  /* fppowbf16.vhdl:1031:23  */
  assign n3685 = x == 10'b0011001001;
  /* fppowbf16.vhdl:1032:23  */
  assign n3688 = x == 10'b0011001010;
  /* fppowbf16.vhdl:1033:23  */
  assign n3691 = x == 10'b0011001011;
  /* fppowbf16.vhdl:1034:23  */
  assign n3694 = x == 10'b0011001100;
  /* fppowbf16.vhdl:1035:23  */
  assign n3697 = x == 10'b0011001101;
  /* fppowbf16.vhdl:1036:23  */
  assign n3700 = x == 10'b0011001110;
  /* fppowbf16.vhdl:1037:23  */
  assign n3703 = x == 10'b0011001111;
  /* fppowbf16.vhdl:1038:23  */
  assign n3706 = x == 10'b0011010000;
  /* fppowbf16.vhdl:1039:23  */
  assign n3709 = x == 10'b0011010001;
  /* fppowbf16.vhdl:1040:23  */
  assign n3712 = x == 10'b0011010010;
  /* fppowbf16.vhdl:1041:23  */
  assign n3715 = x == 10'b0011010011;
  /* fppowbf16.vhdl:1042:23  */
  assign n3718 = x == 10'b0011010100;
  /* fppowbf16.vhdl:1043:23  */
  assign n3721 = x == 10'b0011010101;
  /* fppowbf16.vhdl:1044:23  */
  assign n3724 = x == 10'b0011010110;
  /* fppowbf16.vhdl:1045:23  */
  assign n3727 = x == 10'b0011010111;
  /* fppowbf16.vhdl:1046:23  */
  assign n3730 = x == 10'b0011011000;
  /* fppowbf16.vhdl:1047:23  */
  assign n3733 = x == 10'b0011011001;
  /* fppowbf16.vhdl:1048:23  */
  assign n3736 = x == 10'b0011011010;
  /* fppowbf16.vhdl:1049:23  */
  assign n3739 = x == 10'b0011011011;
  /* fppowbf16.vhdl:1050:23  */
  assign n3742 = x == 10'b0011011100;
  /* fppowbf16.vhdl:1051:23  */
  assign n3745 = x == 10'b0011011101;
  /* fppowbf16.vhdl:1052:23  */
  assign n3748 = x == 10'b0011011110;
  /* fppowbf16.vhdl:1053:23  */
  assign n3751 = x == 10'b0011011111;
  /* fppowbf16.vhdl:1054:23  */
  assign n3754 = x == 10'b0011100000;
  /* fppowbf16.vhdl:1055:23  */
  assign n3757 = x == 10'b0011100001;
  /* fppowbf16.vhdl:1056:23  */
  assign n3760 = x == 10'b0011100010;
  /* fppowbf16.vhdl:1057:23  */
  assign n3763 = x == 10'b0011100011;
  /* fppowbf16.vhdl:1058:23  */
  assign n3766 = x == 10'b0011100100;
  /* fppowbf16.vhdl:1059:23  */
  assign n3769 = x == 10'b0011100101;
  /* fppowbf16.vhdl:1060:23  */
  assign n3772 = x == 10'b0011100110;
  /* fppowbf16.vhdl:1061:23  */
  assign n3775 = x == 10'b0011100111;
  /* fppowbf16.vhdl:1062:23  */
  assign n3778 = x == 10'b0011101000;
  /* fppowbf16.vhdl:1063:23  */
  assign n3781 = x == 10'b0011101001;
  /* fppowbf16.vhdl:1064:23  */
  assign n3784 = x == 10'b0011101010;
  /* fppowbf16.vhdl:1065:23  */
  assign n3787 = x == 10'b0011101011;
  /* fppowbf16.vhdl:1066:23  */
  assign n3790 = x == 10'b0011101100;
  /* fppowbf16.vhdl:1067:23  */
  assign n3793 = x == 10'b0011101101;
  /* fppowbf16.vhdl:1068:23  */
  assign n3796 = x == 10'b0011101110;
  /* fppowbf16.vhdl:1069:23  */
  assign n3799 = x == 10'b0011101111;
  /* fppowbf16.vhdl:1070:23  */
  assign n3802 = x == 10'b0011110000;
  /* fppowbf16.vhdl:1071:23  */
  assign n3805 = x == 10'b0011110001;
  /* fppowbf16.vhdl:1072:23  */
  assign n3808 = x == 10'b0011110010;
  /* fppowbf16.vhdl:1073:23  */
  assign n3811 = x == 10'b0011110011;
  /* fppowbf16.vhdl:1074:23  */
  assign n3814 = x == 10'b0011110100;
  /* fppowbf16.vhdl:1075:23  */
  assign n3817 = x == 10'b0011110101;
  /* fppowbf16.vhdl:1076:23  */
  assign n3820 = x == 10'b0011110110;
  /* fppowbf16.vhdl:1077:23  */
  assign n3823 = x == 10'b0011110111;
  /* fppowbf16.vhdl:1078:23  */
  assign n3826 = x == 10'b0011111000;
  /* fppowbf16.vhdl:1079:23  */
  assign n3829 = x == 10'b0011111001;
  /* fppowbf16.vhdl:1080:23  */
  assign n3832 = x == 10'b0011111010;
  /* fppowbf16.vhdl:1081:23  */
  assign n3835 = x == 10'b0011111011;
  /* fppowbf16.vhdl:1082:23  */
  assign n3838 = x == 10'b0011111100;
  /* fppowbf16.vhdl:1083:23  */
  assign n3841 = x == 10'b0011111101;
  /* fppowbf16.vhdl:1084:23  */
  assign n3844 = x == 10'b0011111110;
  /* fppowbf16.vhdl:1085:23  */
  assign n3847 = x == 10'b0011111111;
  /* fppowbf16.vhdl:1086:23  */
  assign n3850 = x == 10'b0100000000;
  /* fppowbf16.vhdl:1087:23  */
  assign n3853 = x == 10'b0100000001;
  /* fppowbf16.vhdl:1088:23  */
  assign n3856 = x == 10'b0100000010;
  /* fppowbf16.vhdl:1089:23  */
  assign n3859 = x == 10'b0100000011;
  /* fppowbf16.vhdl:1090:23  */
  assign n3862 = x == 10'b0100000100;
  /* fppowbf16.vhdl:1091:23  */
  assign n3865 = x == 10'b0100000101;
  /* fppowbf16.vhdl:1092:23  */
  assign n3868 = x == 10'b0100000110;
  /* fppowbf16.vhdl:1093:23  */
  assign n3871 = x == 10'b0100000111;
  /* fppowbf16.vhdl:1094:23  */
  assign n3874 = x == 10'b0100001000;
  /* fppowbf16.vhdl:1095:23  */
  assign n3877 = x == 10'b0100001001;
  /* fppowbf16.vhdl:1096:23  */
  assign n3880 = x == 10'b0100001010;
  /* fppowbf16.vhdl:1097:23  */
  assign n3883 = x == 10'b0100001011;
  /* fppowbf16.vhdl:1098:23  */
  assign n3886 = x == 10'b0100001100;
  /* fppowbf16.vhdl:1099:23  */
  assign n3889 = x == 10'b0100001101;
  /* fppowbf16.vhdl:1100:23  */
  assign n3892 = x == 10'b0100001110;
  /* fppowbf16.vhdl:1101:23  */
  assign n3895 = x == 10'b0100001111;
  /* fppowbf16.vhdl:1102:23  */
  assign n3898 = x == 10'b0100010000;
  /* fppowbf16.vhdl:1103:23  */
  assign n3901 = x == 10'b0100010001;
  /* fppowbf16.vhdl:1104:23  */
  assign n3904 = x == 10'b0100010010;
  /* fppowbf16.vhdl:1105:23  */
  assign n3907 = x == 10'b0100010011;
  /* fppowbf16.vhdl:1106:23  */
  assign n3910 = x == 10'b0100010100;
  /* fppowbf16.vhdl:1107:23  */
  assign n3913 = x == 10'b0100010101;
  /* fppowbf16.vhdl:1108:23  */
  assign n3916 = x == 10'b0100010110;
  /* fppowbf16.vhdl:1109:23  */
  assign n3919 = x == 10'b0100010111;
  /* fppowbf16.vhdl:1110:23  */
  assign n3922 = x == 10'b0100011000;
  /* fppowbf16.vhdl:1111:23  */
  assign n3925 = x == 10'b0100011001;
  /* fppowbf16.vhdl:1112:23  */
  assign n3928 = x == 10'b0100011010;
  /* fppowbf16.vhdl:1113:23  */
  assign n3931 = x == 10'b0100011011;
  /* fppowbf16.vhdl:1114:23  */
  assign n3934 = x == 10'b0100011100;
  /* fppowbf16.vhdl:1115:23  */
  assign n3937 = x == 10'b0100011101;
  /* fppowbf16.vhdl:1116:23  */
  assign n3940 = x == 10'b0100011110;
  /* fppowbf16.vhdl:1117:23  */
  assign n3943 = x == 10'b0100011111;
  /* fppowbf16.vhdl:1118:23  */
  assign n3946 = x == 10'b0100100000;
  /* fppowbf16.vhdl:1119:23  */
  assign n3949 = x == 10'b0100100001;
  /* fppowbf16.vhdl:1120:23  */
  assign n3952 = x == 10'b0100100010;
  /* fppowbf16.vhdl:1121:23  */
  assign n3955 = x == 10'b0100100011;
  /* fppowbf16.vhdl:1122:23  */
  assign n3958 = x == 10'b0100100100;
  /* fppowbf16.vhdl:1123:23  */
  assign n3961 = x == 10'b0100100101;
  /* fppowbf16.vhdl:1124:23  */
  assign n3964 = x == 10'b0100100110;
  /* fppowbf16.vhdl:1125:23  */
  assign n3967 = x == 10'b0100100111;
  /* fppowbf16.vhdl:1126:23  */
  assign n3970 = x == 10'b0100101000;
  /* fppowbf16.vhdl:1127:23  */
  assign n3973 = x == 10'b0100101001;
  /* fppowbf16.vhdl:1128:23  */
  assign n3976 = x == 10'b0100101010;
  /* fppowbf16.vhdl:1129:23  */
  assign n3979 = x == 10'b0100101011;
  /* fppowbf16.vhdl:1130:23  */
  assign n3982 = x == 10'b0100101100;
  /* fppowbf16.vhdl:1131:23  */
  assign n3985 = x == 10'b0100101101;
  /* fppowbf16.vhdl:1132:23  */
  assign n3988 = x == 10'b0100101110;
  /* fppowbf16.vhdl:1133:23  */
  assign n3991 = x == 10'b0100101111;
  /* fppowbf16.vhdl:1134:23  */
  assign n3994 = x == 10'b0100110000;
  /* fppowbf16.vhdl:1135:23  */
  assign n3997 = x == 10'b0100110001;
  /* fppowbf16.vhdl:1136:23  */
  assign n4000 = x == 10'b0100110010;
  /* fppowbf16.vhdl:1137:23  */
  assign n4003 = x == 10'b0100110011;
  /* fppowbf16.vhdl:1138:23  */
  assign n4006 = x == 10'b0100110100;
  /* fppowbf16.vhdl:1139:23  */
  assign n4009 = x == 10'b0100110101;
  /* fppowbf16.vhdl:1140:23  */
  assign n4012 = x == 10'b0100110110;
  /* fppowbf16.vhdl:1141:23  */
  assign n4015 = x == 10'b0100110111;
  /* fppowbf16.vhdl:1142:23  */
  assign n4018 = x == 10'b0100111000;
  /* fppowbf16.vhdl:1143:23  */
  assign n4021 = x == 10'b0100111001;
  /* fppowbf16.vhdl:1144:23  */
  assign n4024 = x == 10'b0100111010;
  /* fppowbf16.vhdl:1145:23  */
  assign n4027 = x == 10'b0100111011;
  /* fppowbf16.vhdl:1146:23  */
  assign n4030 = x == 10'b0100111100;
  /* fppowbf16.vhdl:1147:23  */
  assign n4033 = x == 10'b0100111101;
  /* fppowbf16.vhdl:1148:23  */
  assign n4036 = x == 10'b0100111110;
  /* fppowbf16.vhdl:1149:23  */
  assign n4039 = x == 10'b0100111111;
  /* fppowbf16.vhdl:1150:23  */
  assign n4042 = x == 10'b0101000000;
  /* fppowbf16.vhdl:1151:23  */
  assign n4045 = x == 10'b0101000001;
  /* fppowbf16.vhdl:1152:23  */
  assign n4048 = x == 10'b0101000010;
  /* fppowbf16.vhdl:1153:23  */
  assign n4051 = x == 10'b0101000011;
  /* fppowbf16.vhdl:1154:23  */
  assign n4054 = x == 10'b0101000100;
  /* fppowbf16.vhdl:1155:23  */
  assign n4057 = x == 10'b0101000101;
  /* fppowbf16.vhdl:1156:23  */
  assign n4060 = x == 10'b0101000110;
  /* fppowbf16.vhdl:1157:23  */
  assign n4063 = x == 10'b0101000111;
  /* fppowbf16.vhdl:1158:23  */
  assign n4066 = x == 10'b0101001000;
  /* fppowbf16.vhdl:1159:23  */
  assign n4069 = x == 10'b0101001001;
  /* fppowbf16.vhdl:1160:23  */
  assign n4072 = x == 10'b0101001010;
  /* fppowbf16.vhdl:1161:23  */
  assign n4075 = x == 10'b0101001011;
  /* fppowbf16.vhdl:1162:23  */
  assign n4078 = x == 10'b0101001100;
  /* fppowbf16.vhdl:1163:23  */
  assign n4081 = x == 10'b0101001101;
  /* fppowbf16.vhdl:1164:23  */
  assign n4084 = x == 10'b0101001110;
  /* fppowbf16.vhdl:1165:23  */
  assign n4087 = x == 10'b0101001111;
  /* fppowbf16.vhdl:1166:23  */
  assign n4090 = x == 10'b0101010000;
  /* fppowbf16.vhdl:1167:23  */
  assign n4093 = x == 10'b0101010001;
  /* fppowbf16.vhdl:1168:23  */
  assign n4096 = x == 10'b0101010010;
  /* fppowbf16.vhdl:1169:23  */
  assign n4099 = x == 10'b0101010011;
  /* fppowbf16.vhdl:1170:23  */
  assign n4102 = x == 10'b0101010100;
  /* fppowbf16.vhdl:1171:23  */
  assign n4105 = x == 10'b0101010101;
  /* fppowbf16.vhdl:1172:23  */
  assign n4108 = x == 10'b0101010110;
  /* fppowbf16.vhdl:1173:23  */
  assign n4111 = x == 10'b0101010111;
  /* fppowbf16.vhdl:1174:23  */
  assign n4114 = x == 10'b0101011000;
  /* fppowbf16.vhdl:1175:23  */
  assign n4117 = x == 10'b0101011001;
  /* fppowbf16.vhdl:1176:23  */
  assign n4120 = x == 10'b0101011010;
  /* fppowbf16.vhdl:1177:23  */
  assign n4123 = x == 10'b0101011011;
  /* fppowbf16.vhdl:1178:23  */
  assign n4126 = x == 10'b0101011100;
  /* fppowbf16.vhdl:1179:23  */
  assign n4129 = x == 10'b0101011101;
  /* fppowbf16.vhdl:1180:23  */
  assign n4132 = x == 10'b0101011110;
  /* fppowbf16.vhdl:1181:23  */
  assign n4135 = x == 10'b0101011111;
  /* fppowbf16.vhdl:1182:23  */
  assign n4138 = x == 10'b0101100000;
  /* fppowbf16.vhdl:1183:23  */
  assign n4141 = x == 10'b0101100001;
  /* fppowbf16.vhdl:1184:23  */
  assign n4144 = x == 10'b0101100010;
  /* fppowbf16.vhdl:1185:23  */
  assign n4147 = x == 10'b0101100011;
  /* fppowbf16.vhdl:1186:23  */
  assign n4150 = x == 10'b0101100100;
  /* fppowbf16.vhdl:1187:23  */
  assign n4153 = x == 10'b0101100101;
  /* fppowbf16.vhdl:1188:23  */
  assign n4156 = x == 10'b0101100110;
  /* fppowbf16.vhdl:1189:23  */
  assign n4159 = x == 10'b0101100111;
  /* fppowbf16.vhdl:1190:23  */
  assign n4162 = x == 10'b0101101000;
  /* fppowbf16.vhdl:1191:23  */
  assign n4165 = x == 10'b0101101001;
  /* fppowbf16.vhdl:1192:23  */
  assign n4168 = x == 10'b0101101010;
  /* fppowbf16.vhdl:1193:23  */
  assign n4171 = x == 10'b0101101011;
  /* fppowbf16.vhdl:1194:23  */
  assign n4174 = x == 10'b0101101100;
  /* fppowbf16.vhdl:1195:23  */
  assign n4177 = x == 10'b0101101101;
  /* fppowbf16.vhdl:1196:23  */
  assign n4180 = x == 10'b0101101110;
  /* fppowbf16.vhdl:1197:23  */
  assign n4183 = x == 10'b0101101111;
  /* fppowbf16.vhdl:1198:23  */
  assign n4186 = x == 10'b0101110000;
  /* fppowbf16.vhdl:1199:23  */
  assign n4189 = x == 10'b0101110001;
  /* fppowbf16.vhdl:1200:23  */
  assign n4192 = x == 10'b0101110010;
  /* fppowbf16.vhdl:1201:23  */
  assign n4195 = x == 10'b0101110011;
  /* fppowbf16.vhdl:1202:23  */
  assign n4198 = x == 10'b0101110100;
  /* fppowbf16.vhdl:1203:23  */
  assign n4201 = x == 10'b0101110101;
  /* fppowbf16.vhdl:1204:23  */
  assign n4204 = x == 10'b0101110110;
  /* fppowbf16.vhdl:1205:23  */
  assign n4207 = x == 10'b0101110111;
  /* fppowbf16.vhdl:1206:23  */
  assign n4210 = x == 10'b0101111000;
  /* fppowbf16.vhdl:1207:23  */
  assign n4213 = x == 10'b0101111001;
  /* fppowbf16.vhdl:1208:23  */
  assign n4216 = x == 10'b0101111010;
  /* fppowbf16.vhdl:1209:23  */
  assign n4219 = x == 10'b0101111011;
  /* fppowbf16.vhdl:1210:23  */
  assign n4222 = x == 10'b0101111100;
  /* fppowbf16.vhdl:1211:23  */
  assign n4225 = x == 10'b0101111101;
  /* fppowbf16.vhdl:1212:23  */
  assign n4228 = x == 10'b0101111110;
  /* fppowbf16.vhdl:1213:23  */
  assign n4231 = x == 10'b0101111111;
  /* fppowbf16.vhdl:1214:23  */
  assign n4234 = x == 10'b0110000000;
  /* fppowbf16.vhdl:1215:23  */
  assign n4237 = x == 10'b0110000001;
  /* fppowbf16.vhdl:1216:23  */
  assign n4240 = x == 10'b0110000010;
  /* fppowbf16.vhdl:1217:23  */
  assign n4243 = x == 10'b0110000011;
  /* fppowbf16.vhdl:1218:23  */
  assign n4246 = x == 10'b0110000100;
  /* fppowbf16.vhdl:1219:23  */
  assign n4249 = x == 10'b0110000101;
  /* fppowbf16.vhdl:1220:23  */
  assign n4252 = x == 10'b0110000110;
  /* fppowbf16.vhdl:1221:23  */
  assign n4255 = x == 10'b0110000111;
  /* fppowbf16.vhdl:1222:23  */
  assign n4258 = x == 10'b0110001000;
  /* fppowbf16.vhdl:1223:23  */
  assign n4261 = x == 10'b0110001001;
  /* fppowbf16.vhdl:1224:23  */
  assign n4264 = x == 10'b0110001010;
  /* fppowbf16.vhdl:1225:23  */
  assign n4267 = x == 10'b0110001011;
  /* fppowbf16.vhdl:1226:23  */
  assign n4270 = x == 10'b0110001100;
  /* fppowbf16.vhdl:1227:23  */
  assign n4273 = x == 10'b0110001101;
  /* fppowbf16.vhdl:1228:23  */
  assign n4276 = x == 10'b0110001110;
  /* fppowbf16.vhdl:1229:23  */
  assign n4279 = x == 10'b0110001111;
  /* fppowbf16.vhdl:1230:23  */
  assign n4282 = x == 10'b0110010000;
  /* fppowbf16.vhdl:1231:23  */
  assign n4285 = x == 10'b0110010001;
  /* fppowbf16.vhdl:1232:23  */
  assign n4288 = x == 10'b0110010010;
  /* fppowbf16.vhdl:1233:23  */
  assign n4291 = x == 10'b0110010011;
  /* fppowbf16.vhdl:1234:23  */
  assign n4294 = x == 10'b0110010100;
  /* fppowbf16.vhdl:1235:23  */
  assign n4297 = x == 10'b0110010101;
  /* fppowbf16.vhdl:1236:23  */
  assign n4300 = x == 10'b0110010110;
  /* fppowbf16.vhdl:1237:23  */
  assign n4303 = x == 10'b0110010111;
  /* fppowbf16.vhdl:1238:23  */
  assign n4306 = x == 10'b0110011000;
  /* fppowbf16.vhdl:1239:23  */
  assign n4309 = x == 10'b0110011001;
  /* fppowbf16.vhdl:1240:23  */
  assign n4312 = x == 10'b0110011010;
  /* fppowbf16.vhdl:1241:23  */
  assign n4315 = x == 10'b0110011011;
  /* fppowbf16.vhdl:1242:23  */
  assign n4318 = x == 10'b0110011100;
  /* fppowbf16.vhdl:1243:23  */
  assign n4321 = x == 10'b0110011101;
  /* fppowbf16.vhdl:1244:23  */
  assign n4324 = x == 10'b0110011110;
  /* fppowbf16.vhdl:1245:23  */
  assign n4327 = x == 10'b0110011111;
  /* fppowbf16.vhdl:1246:23  */
  assign n4330 = x == 10'b0110100000;
  /* fppowbf16.vhdl:1247:23  */
  assign n4333 = x == 10'b0110100001;
  /* fppowbf16.vhdl:1248:23  */
  assign n4336 = x == 10'b0110100010;
  /* fppowbf16.vhdl:1249:23  */
  assign n4339 = x == 10'b0110100011;
  /* fppowbf16.vhdl:1250:23  */
  assign n4342 = x == 10'b0110100100;
  /* fppowbf16.vhdl:1251:23  */
  assign n4345 = x == 10'b0110100101;
  /* fppowbf16.vhdl:1252:23  */
  assign n4348 = x == 10'b0110100110;
  /* fppowbf16.vhdl:1253:23  */
  assign n4351 = x == 10'b0110100111;
  /* fppowbf16.vhdl:1254:23  */
  assign n4354 = x == 10'b0110101000;
  /* fppowbf16.vhdl:1255:23  */
  assign n4357 = x == 10'b0110101001;
  /* fppowbf16.vhdl:1256:23  */
  assign n4360 = x == 10'b0110101010;
  /* fppowbf16.vhdl:1257:23  */
  assign n4363 = x == 10'b0110101011;
  /* fppowbf16.vhdl:1258:23  */
  assign n4366 = x == 10'b0110101100;
  /* fppowbf16.vhdl:1259:23  */
  assign n4369 = x == 10'b0110101101;
  /* fppowbf16.vhdl:1260:23  */
  assign n4372 = x == 10'b0110101110;
  /* fppowbf16.vhdl:1261:23  */
  assign n4375 = x == 10'b0110101111;
  /* fppowbf16.vhdl:1262:23  */
  assign n4378 = x == 10'b0110110000;
  /* fppowbf16.vhdl:1263:23  */
  assign n4381 = x == 10'b0110110001;
  /* fppowbf16.vhdl:1264:23  */
  assign n4384 = x == 10'b0110110010;
  /* fppowbf16.vhdl:1265:23  */
  assign n4387 = x == 10'b0110110011;
  /* fppowbf16.vhdl:1266:23  */
  assign n4390 = x == 10'b0110110100;
  /* fppowbf16.vhdl:1267:23  */
  assign n4393 = x == 10'b0110110101;
  /* fppowbf16.vhdl:1268:23  */
  assign n4396 = x == 10'b0110110110;
  /* fppowbf16.vhdl:1269:23  */
  assign n4399 = x == 10'b0110110111;
  /* fppowbf16.vhdl:1270:23  */
  assign n4402 = x == 10'b0110111000;
  /* fppowbf16.vhdl:1271:23  */
  assign n4405 = x == 10'b0110111001;
  /* fppowbf16.vhdl:1272:23  */
  assign n4408 = x == 10'b0110111010;
  /* fppowbf16.vhdl:1273:23  */
  assign n4411 = x == 10'b0110111011;
  /* fppowbf16.vhdl:1274:23  */
  assign n4414 = x == 10'b0110111100;
  /* fppowbf16.vhdl:1275:23  */
  assign n4417 = x == 10'b0110111101;
  /* fppowbf16.vhdl:1276:23  */
  assign n4420 = x == 10'b0110111110;
  /* fppowbf16.vhdl:1277:23  */
  assign n4423 = x == 10'b0110111111;
  /* fppowbf16.vhdl:1278:23  */
  assign n4426 = x == 10'b0111000000;
  /* fppowbf16.vhdl:1279:23  */
  assign n4429 = x == 10'b0111000001;
  /* fppowbf16.vhdl:1280:23  */
  assign n4432 = x == 10'b0111000010;
  /* fppowbf16.vhdl:1281:23  */
  assign n4435 = x == 10'b0111000011;
  /* fppowbf16.vhdl:1282:23  */
  assign n4438 = x == 10'b0111000100;
  /* fppowbf16.vhdl:1283:23  */
  assign n4441 = x == 10'b0111000101;
  /* fppowbf16.vhdl:1284:23  */
  assign n4444 = x == 10'b0111000110;
  /* fppowbf16.vhdl:1285:23  */
  assign n4447 = x == 10'b0111000111;
  /* fppowbf16.vhdl:1286:23  */
  assign n4450 = x == 10'b0111001000;
  /* fppowbf16.vhdl:1287:23  */
  assign n4453 = x == 10'b0111001001;
  /* fppowbf16.vhdl:1288:23  */
  assign n4456 = x == 10'b0111001010;
  /* fppowbf16.vhdl:1289:23  */
  assign n4459 = x == 10'b0111001011;
  /* fppowbf16.vhdl:1290:23  */
  assign n4462 = x == 10'b0111001100;
  /* fppowbf16.vhdl:1291:23  */
  assign n4465 = x == 10'b0111001101;
  /* fppowbf16.vhdl:1292:23  */
  assign n4468 = x == 10'b0111001110;
  /* fppowbf16.vhdl:1293:23  */
  assign n4471 = x == 10'b0111001111;
  /* fppowbf16.vhdl:1294:23  */
  assign n4474 = x == 10'b0111010000;
  /* fppowbf16.vhdl:1295:23  */
  assign n4477 = x == 10'b0111010001;
  /* fppowbf16.vhdl:1296:23  */
  assign n4480 = x == 10'b0111010010;
  /* fppowbf16.vhdl:1297:23  */
  assign n4483 = x == 10'b0111010011;
  /* fppowbf16.vhdl:1298:23  */
  assign n4486 = x == 10'b0111010100;
  /* fppowbf16.vhdl:1299:23  */
  assign n4489 = x == 10'b0111010101;
  /* fppowbf16.vhdl:1300:23  */
  assign n4492 = x == 10'b0111010110;
  /* fppowbf16.vhdl:1301:23  */
  assign n4495 = x == 10'b0111010111;
  /* fppowbf16.vhdl:1302:23  */
  assign n4498 = x == 10'b0111011000;
  /* fppowbf16.vhdl:1303:23  */
  assign n4501 = x == 10'b0111011001;
  /* fppowbf16.vhdl:1304:23  */
  assign n4504 = x == 10'b0111011010;
  /* fppowbf16.vhdl:1305:23  */
  assign n4507 = x == 10'b0111011011;
  /* fppowbf16.vhdl:1306:23  */
  assign n4510 = x == 10'b0111011100;
  /* fppowbf16.vhdl:1307:23  */
  assign n4513 = x == 10'b0111011101;
  /* fppowbf16.vhdl:1308:23  */
  assign n4516 = x == 10'b0111011110;
  /* fppowbf16.vhdl:1309:23  */
  assign n4519 = x == 10'b0111011111;
  /* fppowbf16.vhdl:1310:23  */
  assign n4522 = x == 10'b0111100000;
  /* fppowbf16.vhdl:1311:23  */
  assign n4525 = x == 10'b0111100001;
  /* fppowbf16.vhdl:1312:23  */
  assign n4528 = x == 10'b0111100010;
  /* fppowbf16.vhdl:1313:23  */
  assign n4531 = x == 10'b0111100011;
  /* fppowbf16.vhdl:1314:23  */
  assign n4534 = x == 10'b0111100100;
  /* fppowbf16.vhdl:1315:23  */
  assign n4537 = x == 10'b0111100101;
  /* fppowbf16.vhdl:1316:23  */
  assign n4540 = x == 10'b0111100110;
  /* fppowbf16.vhdl:1317:23  */
  assign n4543 = x == 10'b0111100111;
  /* fppowbf16.vhdl:1318:23  */
  assign n4546 = x == 10'b0111101000;
  /* fppowbf16.vhdl:1319:23  */
  assign n4549 = x == 10'b0111101001;
  /* fppowbf16.vhdl:1320:23  */
  assign n4552 = x == 10'b0111101010;
  /* fppowbf16.vhdl:1321:23  */
  assign n4555 = x == 10'b0111101011;
  /* fppowbf16.vhdl:1322:23  */
  assign n4558 = x == 10'b0111101100;
  /* fppowbf16.vhdl:1323:23  */
  assign n4561 = x == 10'b0111101101;
  /* fppowbf16.vhdl:1324:23  */
  assign n4564 = x == 10'b0111101110;
  /* fppowbf16.vhdl:1325:23  */
  assign n4567 = x == 10'b0111101111;
  /* fppowbf16.vhdl:1326:23  */
  assign n4570 = x == 10'b0111110000;
  /* fppowbf16.vhdl:1327:23  */
  assign n4573 = x == 10'b0111110001;
  /* fppowbf16.vhdl:1328:23  */
  assign n4576 = x == 10'b0111110010;
  /* fppowbf16.vhdl:1329:23  */
  assign n4579 = x == 10'b0111110011;
  /* fppowbf16.vhdl:1330:23  */
  assign n4582 = x == 10'b0111110100;
  /* fppowbf16.vhdl:1331:23  */
  assign n4585 = x == 10'b0111110101;
  /* fppowbf16.vhdl:1332:23  */
  assign n4588 = x == 10'b0111110110;
  /* fppowbf16.vhdl:1333:23  */
  assign n4591 = x == 10'b0111110111;
  /* fppowbf16.vhdl:1334:23  */
  assign n4594 = x == 10'b0111111000;
  /* fppowbf16.vhdl:1335:23  */
  assign n4597 = x == 10'b0111111001;
  /* fppowbf16.vhdl:1336:23  */
  assign n4600 = x == 10'b0111111010;
  /* fppowbf16.vhdl:1337:23  */
  assign n4603 = x == 10'b0111111011;
  /* fppowbf16.vhdl:1338:23  */
  assign n4606 = x == 10'b0111111100;
  /* fppowbf16.vhdl:1339:23  */
  assign n4609 = x == 10'b0111111101;
  /* fppowbf16.vhdl:1340:23  */
  assign n4612 = x == 10'b0111111110;
  /* fppowbf16.vhdl:1341:23  */
  assign n4615 = x == 10'b0111111111;
  /* fppowbf16.vhdl:1342:23  */
  assign n4618 = x == 10'b1000000000;
  /* fppowbf16.vhdl:1343:23  */
  assign n4621 = x == 10'b1000000001;
  /* fppowbf16.vhdl:1344:23  */
  assign n4624 = x == 10'b1000000010;
  /* fppowbf16.vhdl:1345:23  */
  assign n4627 = x == 10'b1000000011;
  /* fppowbf16.vhdl:1346:23  */
  assign n4630 = x == 10'b1000000100;
  /* fppowbf16.vhdl:1347:23  */
  assign n4633 = x == 10'b1000000101;
  /* fppowbf16.vhdl:1348:23  */
  assign n4636 = x == 10'b1000000110;
  /* fppowbf16.vhdl:1349:23  */
  assign n4639 = x == 10'b1000000111;
  /* fppowbf16.vhdl:1350:23  */
  assign n4642 = x == 10'b1000001000;
  /* fppowbf16.vhdl:1351:23  */
  assign n4645 = x == 10'b1000001001;
  /* fppowbf16.vhdl:1352:23  */
  assign n4648 = x == 10'b1000001010;
  /* fppowbf16.vhdl:1353:23  */
  assign n4651 = x == 10'b1000001011;
  /* fppowbf16.vhdl:1354:23  */
  assign n4654 = x == 10'b1000001100;
  /* fppowbf16.vhdl:1355:23  */
  assign n4657 = x == 10'b1000001101;
  /* fppowbf16.vhdl:1356:23  */
  assign n4660 = x == 10'b1000001110;
  /* fppowbf16.vhdl:1357:23  */
  assign n4663 = x == 10'b1000001111;
  /* fppowbf16.vhdl:1358:23  */
  assign n4666 = x == 10'b1000010000;
  /* fppowbf16.vhdl:1359:23  */
  assign n4669 = x == 10'b1000010001;
  /* fppowbf16.vhdl:1360:23  */
  assign n4672 = x == 10'b1000010010;
  /* fppowbf16.vhdl:1361:23  */
  assign n4675 = x == 10'b1000010011;
  /* fppowbf16.vhdl:1362:23  */
  assign n4678 = x == 10'b1000010100;
  /* fppowbf16.vhdl:1363:23  */
  assign n4681 = x == 10'b1000010101;
  /* fppowbf16.vhdl:1364:23  */
  assign n4684 = x == 10'b1000010110;
  /* fppowbf16.vhdl:1365:23  */
  assign n4687 = x == 10'b1000010111;
  /* fppowbf16.vhdl:1366:23  */
  assign n4690 = x == 10'b1000011000;
  /* fppowbf16.vhdl:1367:23  */
  assign n4693 = x == 10'b1000011001;
  /* fppowbf16.vhdl:1368:23  */
  assign n4696 = x == 10'b1000011010;
  /* fppowbf16.vhdl:1369:23  */
  assign n4699 = x == 10'b1000011011;
  /* fppowbf16.vhdl:1370:23  */
  assign n4702 = x == 10'b1000011100;
  /* fppowbf16.vhdl:1371:23  */
  assign n4705 = x == 10'b1000011101;
  /* fppowbf16.vhdl:1372:23  */
  assign n4708 = x == 10'b1000011110;
  /* fppowbf16.vhdl:1373:23  */
  assign n4711 = x == 10'b1000011111;
  /* fppowbf16.vhdl:1374:23  */
  assign n4714 = x == 10'b1000100000;
  /* fppowbf16.vhdl:1375:23  */
  assign n4717 = x == 10'b1000100001;
  /* fppowbf16.vhdl:1376:23  */
  assign n4720 = x == 10'b1000100010;
  /* fppowbf16.vhdl:1377:23  */
  assign n4723 = x == 10'b1000100011;
  /* fppowbf16.vhdl:1378:23  */
  assign n4726 = x == 10'b1000100100;
  /* fppowbf16.vhdl:1379:23  */
  assign n4729 = x == 10'b1000100101;
  /* fppowbf16.vhdl:1380:23  */
  assign n4732 = x == 10'b1000100110;
  /* fppowbf16.vhdl:1381:23  */
  assign n4735 = x == 10'b1000100111;
  /* fppowbf16.vhdl:1382:23  */
  assign n4738 = x == 10'b1000101000;
  /* fppowbf16.vhdl:1383:23  */
  assign n4741 = x == 10'b1000101001;
  /* fppowbf16.vhdl:1384:23  */
  assign n4744 = x == 10'b1000101010;
  /* fppowbf16.vhdl:1385:23  */
  assign n4747 = x == 10'b1000101011;
  /* fppowbf16.vhdl:1386:23  */
  assign n4750 = x == 10'b1000101100;
  /* fppowbf16.vhdl:1387:23  */
  assign n4753 = x == 10'b1000101101;
  /* fppowbf16.vhdl:1388:23  */
  assign n4756 = x == 10'b1000101110;
  /* fppowbf16.vhdl:1389:23  */
  assign n4759 = x == 10'b1000101111;
  /* fppowbf16.vhdl:1390:23  */
  assign n4762 = x == 10'b1000110000;
  /* fppowbf16.vhdl:1391:23  */
  assign n4765 = x == 10'b1000110001;
  /* fppowbf16.vhdl:1392:23  */
  assign n4768 = x == 10'b1000110010;
  /* fppowbf16.vhdl:1393:23  */
  assign n4771 = x == 10'b1000110011;
  /* fppowbf16.vhdl:1394:23  */
  assign n4774 = x == 10'b1000110100;
  /* fppowbf16.vhdl:1395:23  */
  assign n4777 = x == 10'b1000110101;
  /* fppowbf16.vhdl:1396:23  */
  assign n4780 = x == 10'b1000110110;
  /* fppowbf16.vhdl:1397:23  */
  assign n4783 = x == 10'b1000110111;
  /* fppowbf16.vhdl:1398:23  */
  assign n4786 = x == 10'b1000111000;
  /* fppowbf16.vhdl:1399:23  */
  assign n4789 = x == 10'b1000111001;
  /* fppowbf16.vhdl:1400:23  */
  assign n4792 = x == 10'b1000111010;
  /* fppowbf16.vhdl:1401:23  */
  assign n4795 = x == 10'b1000111011;
  /* fppowbf16.vhdl:1402:23  */
  assign n4798 = x == 10'b1000111100;
  /* fppowbf16.vhdl:1403:23  */
  assign n4801 = x == 10'b1000111101;
  /* fppowbf16.vhdl:1404:23  */
  assign n4804 = x == 10'b1000111110;
  /* fppowbf16.vhdl:1405:23  */
  assign n4807 = x == 10'b1000111111;
  /* fppowbf16.vhdl:1406:23  */
  assign n4810 = x == 10'b1001000000;
  /* fppowbf16.vhdl:1407:23  */
  assign n4813 = x == 10'b1001000001;
  /* fppowbf16.vhdl:1408:23  */
  assign n4816 = x == 10'b1001000010;
  /* fppowbf16.vhdl:1409:23  */
  assign n4819 = x == 10'b1001000011;
  /* fppowbf16.vhdl:1410:23  */
  assign n4822 = x == 10'b1001000100;
  /* fppowbf16.vhdl:1411:23  */
  assign n4825 = x == 10'b1001000101;
  /* fppowbf16.vhdl:1412:23  */
  assign n4828 = x == 10'b1001000110;
  /* fppowbf16.vhdl:1413:23  */
  assign n4831 = x == 10'b1001000111;
  /* fppowbf16.vhdl:1414:23  */
  assign n4834 = x == 10'b1001001000;
  /* fppowbf16.vhdl:1415:23  */
  assign n4837 = x == 10'b1001001001;
  /* fppowbf16.vhdl:1416:23  */
  assign n4840 = x == 10'b1001001010;
  /* fppowbf16.vhdl:1417:23  */
  assign n4843 = x == 10'b1001001011;
  /* fppowbf16.vhdl:1418:23  */
  assign n4846 = x == 10'b1001001100;
  /* fppowbf16.vhdl:1419:23  */
  assign n4849 = x == 10'b1001001101;
  /* fppowbf16.vhdl:1420:23  */
  assign n4852 = x == 10'b1001001110;
  /* fppowbf16.vhdl:1421:23  */
  assign n4855 = x == 10'b1001001111;
  /* fppowbf16.vhdl:1422:23  */
  assign n4858 = x == 10'b1001010000;
  /* fppowbf16.vhdl:1423:23  */
  assign n4861 = x == 10'b1001010001;
  /* fppowbf16.vhdl:1424:23  */
  assign n4864 = x == 10'b1001010010;
  /* fppowbf16.vhdl:1425:23  */
  assign n4867 = x == 10'b1001010011;
  /* fppowbf16.vhdl:1426:23  */
  assign n4870 = x == 10'b1001010100;
  /* fppowbf16.vhdl:1427:23  */
  assign n4873 = x == 10'b1001010101;
  /* fppowbf16.vhdl:1428:23  */
  assign n4876 = x == 10'b1001010110;
  /* fppowbf16.vhdl:1429:23  */
  assign n4879 = x == 10'b1001010111;
  /* fppowbf16.vhdl:1430:23  */
  assign n4882 = x == 10'b1001011000;
  /* fppowbf16.vhdl:1431:23  */
  assign n4885 = x == 10'b1001011001;
  /* fppowbf16.vhdl:1432:23  */
  assign n4888 = x == 10'b1001011010;
  /* fppowbf16.vhdl:1433:23  */
  assign n4891 = x == 10'b1001011011;
  /* fppowbf16.vhdl:1434:23  */
  assign n4894 = x == 10'b1001011100;
  /* fppowbf16.vhdl:1435:23  */
  assign n4897 = x == 10'b1001011101;
  /* fppowbf16.vhdl:1436:23  */
  assign n4900 = x == 10'b1001011110;
  /* fppowbf16.vhdl:1437:23  */
  assign n4903 = x == 10'b1001011111;
  /* fppowbf16.vhdl:1438:23  */
  assign n4906 = x == 10'b1001100000;
  /* fppowbf16.vhdl:1439:23  */
  assign n4909 = x == 10'b1001100001;
  /* fppowbf16.vhdl:1440:23  */
  assign n4912 = x == 10'b1001100010;
  /* fppowbf16.vhdl:1441:23  */
  assign n4915 = x == 10'b1001100011;
  /* fppowbf16.vhdl:1442:23  */
  assign n4918 = x == 10'b1001100100;
  /* fppowbf16.vhdl:1443:23  */
  assign n4921 = x == 10'b1001100101;
  /* fppowbf16.vhdl:1444:23  */
  assign n4924 = x == 10'b1001100110;
  /* fppowbf16.vhdl:1445:23  */
  assign n4927 = x == 10'b1001100111;
  /* fppowbf16.vhdl:1446:23  */
  assign n4930 = x == 10'b1001101000;
  /* fppowbf16.vhdl:1447:23  */
  assign n4933 = x == 10'b1001101001;
  /* fppowbf16.vhdl:1448:23  */
  assign n4936 = x == 10'b1001101010;
  /* fppowbf16.vhdl:1449:23  */
  assign n4939 = x == 10'b1001101011;
  /* fppowbf16.vhdl:1450:23  */
  assign n4942 = x == 10'b1001101100;
  /* fppowbf16.vhdl:1451:23  */
  assign n4945 = x == 10'b1001101101;
  /* fppowbf16.vhdl:1452:23  */
  assign n4948 = x == 10'b1001101110;
  /* fppowbf16.vhdl:1453:23  */
  assign n4951 = x == 10'b1001101111;
  /* fppowbf16.vhdl:1454:23  */
  assign n4954 = x == 10'b1001110000;
  /* fppowbf16.vhdl:1455:23  */
  assign n4957 = x == 10'b1001110001;
  /* fppowbf16.vhdl:1456:23  */
  assign n4960 = x == 10'b1001110010;
  /* fppowbf16.vhdl:1457:23  */
  assign n4963 = x == 10'b1001110011;
  /* fppowbf16.vhdl:1458:23  */
  assign n4966 = x == 10'b1001110100;
  /* fppowbf16.vhdl:1459:23  */
  assign n4969 = x == 10'b1001110101;
  /* fppowbf16.vhdl:1460:23  */
  assign n4972 = x == 10'b1001110110;
  /* fppowbf16.vhdl:1461:23  */
  assign n4975 = x == 10'b1001110111;
  /* fppowbf16.vhdl:1462:23  */
  assign n4978 = x == 10'b1001111000;
  /* fppowbf16.vhdl:1463:23  */
  assign n4981 = x == 10'b1001111001;
  /* fppowbf16.vhdl:1464:23  */
  assign n4984 = x == 10'b1001111010;
  /* fppowbf16.vhdl:1465:23  */
  assign n4987 = x == 10'b1001111011;
  /* fppowbf16.vhdl:1466:23  */
  assign n4990 = x == 10'b1001111100;
  /* fppowbf16.vhdl:1467:23  */
  assign n4993 = x == 10'b1001111101;
  /* fppowbf16.vhdl:1468:23  */
  assign n4996 = x == 10'b1001111110;
  /* fppowbf16.vhdl:1469:23  */
  assign n4999 = x == 10'b1001111111;
  /* fppowbf16.vhdl:1470:23  */
  assign n5002 = x == 10'b1010000000;
  /* fppowbf16.vhdl:1471:23  */
  assign n5005 = x == 10'b1010000001;
  /* fppowbf16.vhdl:1472:23  */
  assign n5008 = x == 10'b1010000010;
  /* fppowbf16.vhdl:1473:23  */
  assign n5011 = x == 10'b1010000011;
  /* fppowbf16.vhdl:1474:23  */
  assign n5014 = x == 10'b1010000100;
  /* fppowbf16.vhdl:1475:23  */
  assign n5017 = x == 10'b1010000101;
  /* fppowbf16.vhdl:1476:23  */
  assign n5020 = x == 10'b1010000110;
  /* fppowbf16.vhdl:1477:23  */
  assign n5023 = x == 10'b1010000111;
  /* fppowbf16.vhdl:1478:23  */
  assign n5026 = x == 10'b1010001000;
  /* fppowbf16.vhdl:1479:23  */
  assign n5029 = x == 10'b1010001001;
  /* fppowbf16.vhdl:1480:23  */
  assign n5032 = x == 10'b1010001010;
  /* fppowbf16.vhdl:1481:23  */
  assign n5035 = x == 10'b1010001011;
  /* fppowbf16.vhdl:1482:23  */
  assign n5038 = x == 10'b1010001100;
  /* fppowbf16.vhdl:1483:23  */
  assign n5041 = x == 10'b1010001101;
  /* fppowbf16.vhdl:1484:23  */
  assign n5044 = x == 10'b1010001110;
  /* fppowbf16.vhdl:1485:23  */
  assign n5047 = x == 10'b1010001111;
  /* fppowbf16.vhdl:1486:23  */
  assign n5050 = x == 10'b1010010000;
  /* fppowbf16.vhdl:1487:23  */
  assign n5053 = x == 10'b1010010001;
  /* fppowbf16.vhdl:1488:23  */
  assign n5056 = x == 10'b1010010010;
  /* fppowbf16.vhdl:1489:23  */
  assign n5059 = x == 10'b1010010011;
  /* fppowbf16.vhdl:1490:23  */
  assign n5062 = x == 10'b1010010100;
  /* fppowbf16.vhdl:1491:23  */
  assign n5065 = x == 10'b1010010101;
  /* fppowbf16.vhdl:1492:23  */
  assign n5068 = x == 10'b1010010110;
  /* fppowbf16.vhdl:1493:23  */
  assign n5071 = x == 10'b1010010111;
  /* fppowbf16.vhdl:1494:23  */
  assign n5074 = x == 10'b1010011000;
  /* fppowbf16.vhdl:1495:23  */
  assign n5077 = x == 10'b1010011001;
  /* fppowbf16.vhdl:1496:23  */
  assign n5080 = x == 10'b1010011010;
  /* fppowbf16.vhdl:1497:23  */
  assign n5083 = x == 10'b1010011011;
  /* fppowbf16.vhdl:1498:23  */
  assign n5086 = x == 10'b1010011100;
  /* fppowbf16.vhdl:1499:23  */
  assign n5089 = x == 10'b1010011101;
  /* fppowbf16.vhdl:1500:23  */
  assign n5092 = x == 10'b1010011110;
  /* fppowbf16.vhdl:1501:23  */
  assign n5095 = x == 10'b1010011111;
  /* fppowbf16.vhdl:1502:23  */
  assign n5098 = x == 10'b1010100000;
  /* fppowbf16.vhdl:1503:23  */
  assign n5101 = x == 10'b1010100001;
  /* fppowbf16.vhdl:1504:23  */
  assign n5104 = x == 10'b1010100010;
  /* fppowbf16.vhdl:1505:23  */
  assign n5107 = x == 10'b1010100011;
  /* fppowbf16.vhdl:1506:23  */
  assign n5110 = x == 10'b1010100100;
  /* fppowbf16.vhdl:1507:23  */
  assign n5113 = x == 10'b1010100101;
  /* fppowbf16.vhdl:1508:23  */
  assign n5116 = x == 10'b1010100110;
  /* fppowbf16.vhdl:1509:23  */
  assign n5119 = x == 10'b1010100111;
  /* fppowbf16.vhdl:1510:23  */
  assign n5122 = x == 10'b1010101000;
  /* fppowbf16.vhdl:1511:23  */
  assign n5125 = x == 10'b1010101001;
  /* fppowbf16.vhdl:1512:23  */
  assign n5128 = x == 10'b1010101010;
  /* fppowbf16.vhdl:1513:23  */
  assign n5131 = x == 10'b1010101011;
  /* fppowbf16.vhdl:1514:23  */
  assign n5134 = x == 10'b1010101100;
  /* fppowbf16.vhdl:1515:23  */
  assign n5137 = x == 10'b1010101101;
  /* fppowbf16.vhdl:1516:23  */
  assign n5140 = x == 10'b1010101110;
  /* fppowbf16.vhdl:1517:23  */
  assign n5143 = x == 10'b1010101111;
  /* fppowbf16.vhdl:1518:23  */
  assign n5146 = x == 10'b1010110000;
  /* fppowbf16.vhdl:1519:23  */
  assign n5149 = x == 10'b1010110001;
  /* fppowbf16.vhdl:1520:23  */
  assign n5152 = x == 10'b1010110010;
  /* fppowbf16.vhdl:1521:23  */
  assign n5155 = x == 10'b1010110011;
  /* fppowbf16.vhdl:1522:23  */
  assign n5158 = x == 10'b1010110100;
  /* fppowbf16.vhdl:1523:23  */
  assign n5161 = x == 10'b1010110101;
  /* fppowbf16.vhdl:1524:23  */
  assign n5164 = x == 10'b1010110110;
  /* fppowbf16.vhdl:1525:23  */
  assign n5167 = x == 10'b1010110111;
  /* fppowbf16.vhdl:1526:23  */
  assign n5170 = x == 10'b1010111000;
  /* fppowbf16.vhdl:1527:23  */
  assign n5173 = x == 10'b1010111001;
  /* fppowbf16.vhdl:1528:23  */
  assign n5176 = x == 10'b1010111010;
  /* fppowbf16.vhdl:1529:23  */
  assign n5179 = x == 10'b1010111011;
  /* fppowbf16.vhdl:1530:23  */
  assign n5182 = x == 10'b1010111100;
  /* fppowbf16.vhdl:1531:23  */
  assign n5185 = x == 10'b1010111101;
  /* fppowbf16.vhdl:1532:23  */
  assign n5188 = x == 10'b1010111110;
  /* fppowbf16.vhdl:1533:23  */
  assign n5191 = x == 10'b1010111111;
  /* fppowbf16.vhdl:1534:23  */
  assign n5194 = x == 10'b1011000000;
  /* fppowbf16.vhdl:1535:23  */
  assign n5197 = x == 10'b1011000001;
  /* fppowbf16.vhdl:1536:23  */
  assign n5200 = x == 10'b1011000010;
  /* fppowbf16.vhdl:1537:23  */
  assign n5203 = x == 10'b1011000011;
  /* fppowbf16.vhdl:1538:23  */
  assign n5206 = x == 10'b1011000100;
  /* fppowbf16.vhdl:1539:23  */
  assign n5209 = x == 10'b1011000101;
  /* fppowbf16.vhdl:1540:23  */
  assign n5212 = x == 10'b1011000110;
  /* fppowbf16.vhdl:1541:23  */
  assign n5215 = x == 10'b1011000111;
  /* fppowbf16.vhdl:1542:23  */
  assign n5218 = x == 10'b1011001000;
  /* fppowbf16.vhdl:1543:23  */
  assign n5221 = x == 10'b1011001001;
  /* fppowbf16.vhdl:1544:23  */
  assign n5224 = x == 10'b1011001010;
  /* fppowbf16.vhdl:1545:23  */
  assign n5227 = x == 10'b1011001011;
  /* fppowbf16.vhdl:1546:23  */
  assign n5230 = x == 10'b1011001100;
  /* fppowbf16.vhdl:1547:23  */
  assign n5233 = x == 10'b1011001101;
  /* fppowbf16.vhdl:1548:23  */
  assign n5236 = x == 10'b1011001110;
  /* fppowbf16.vhdl:1549:23  */
  assign n5239 = x == 10'b1011001111;
  /* fppowbf16.vhdl:1550:23  */
  assign n5242 = x == 10'b1011010000;
  /* fppowbf16.vhdl:1551:23  */
  assign n5245 = x == 10'b1011010001;
  /* fppowbf16.vhdl:1552:23  */
  assign n5248 = x == 10'b1011010010;
  /* fppowbf16.vhdl:1553:23  */
  assign n5251 = x == 10'b1011010011;
  /* fppowbf16.vhdl:1554:23  */
  assign n5254 = x == 10'b1011010100;
  /* fppowbf16.vhdl:1555:23  */
  assign n5257 = x == 10'b1011010101;
  /* fppowbf16.vhdl:1556:23  */
  assign n5260 = x == 10'b1011010110;
  /* fppowbf16.vhdl:1557:23  */
  assign n5263 = x == 10'b1011010111;
  /* fppowbf16.vhdl:1558:23  */
  assign n5266 = x == 10'b1011011000;
  /* fppowbf16.vhdl:1559:23  */
  assign n5269 = x == 10'b1011011001;
  /* fppowbf16.vhdl:1560:23  */
  assign n5272 = x == 10'b1011011010;
  /* fppowbf16.vhdl:1561:23  */
  assign n5275 = x == 10'b1011011011;
  /* fppowbf16.vhdl:1562:23  */
  assign n5278 = x == 10'b1011011100;
  /* fppowbf16.vhdl:1563:23  */
  assign n5281 = x == 10'b1011011101;
  /* fppowbf16.vhdl:1564:23  */
  assign n5284 = x == 10'b1011011110;
  /* fppowbf16.vhdl:1565:23  */
  assign n5287 = x == 10'b1011011111;
  /* fppowbf16.vhdl:1566:23  */
  assign n5290 = x == 10'b1011100000;
  /* fppowbf16.vhdl:1567:23  */
  assign n5293 = x == 10'b1011100001;
  /* fppowbf16.vhdl:1568:23  */
  assign n5296 = x == 10'b1011100010;
  /* fppowbf16.vhdl:1569:23  */
  assign n5299 = x == 10'b1011100011;
  /* fppowbf16.vhdl:1570:23  */
  assign n5302 = x == 10'b1011100100;
  /* fppowbf16.vhdl:1571:23  */
  assign n5305 = x == 10'b1011100101;
  /* fppowbf16.vhdl:1572:23  */
  assign n5308 = x == 10'b1011100110;
  /* fppowbf16.vhdl:1573:23  */
  assign n5311 = x == 10'b1011100111;
  /* fppowbf16.vhdl:1574:23  */
  assign n5314 = x == 10'b1011101000;
  /* fppowbf16.vhdl:1575:23  */
  assign n5317 = x == 10'b1011101001;
  /* fppowbf16.vhdl:1576:23  */
  assign n5320 = x == 10'b1011101010;
  /* fppowbf16.vhdl:1577:23  */
  assign n5323 = x == 10'b1011101011;
  /* fppowbf16.vhdl:1578:23  */
  assign n5326 = x == 10'b1011101100;
  /* fppowbf16.vhdl:1579:23  */
  assign n5329 = x == 10'b1011101101;
  /* fppowbf16.vhdl:1580:23  */
  assign n5332 = x == 10'b1011101110;
  /* fppowbf16.vhdl:1581:23  */
  assign n5335 = x == 10'b1011101111;
  /* fppowbf16.vhdl:1582:23  */
  assign n5338 = x == 10'b1011110000;
  /* fppowbf16.vhdl:1583:23  */
  assign n5341 = x == 10'b1011110001;
  /* fppowbf16.vhdl:1584:23  */
  assign n5344 = x == 10'b1011110010;
  /* fppowbf16.vhdl:1585:23  */
  assign n5347 = x == 10'b1011110011;
  /* fppowbf16.vhdl:1586:23  */
  assign n5350 = x == 10'b1011110100;
  /* fppowbf16.vhdl:1587:23  */
  assign n5353 = x == 10'b1011110101;
  /* fppowbf16.vhdl:1588:23  */
  assign n5356 = x == 10'b1011110110;
  /* fppowbf16.vhdl:1589:23  */
  assign n5359 = x == 10'b1011110111;
  /* fppowbf16.vhdl:1590:23  */
  assign n5362 = x == 10'b1011111000;
  /* fppowbf16.vhdl:1591:23  */
  assign n5365 = x == 10'b1011111001;
  /* fppowbf16.vhdl:1592:23  */
  assign n5368 = x == 10'b1011111010;
  /* fppowbf16.vhdl:1593:23  */
  assign n5371 = x == 10'b1011111011;
  /* fppowbf16.vhdl:1594:23  */
  assign n5374 = x == 10'b1011111100;
  /* fppowbf16.vhdl:1595:23  */
  assign n5377 = x == 10'b1011111101;
  /* fppowbf16.vhdl:1596:23  */
  assign n5380 = x == 10'b1011111110;
  /* fppowbf16.vhdl:1597:23  */
  assign n5383 = x == 10'b1011111111;
  /* fppowbf16.vhdl:1598:23  */
  assign n5386 = x == 10'b1100000000;
  /* fppowbf16.vhdl:1599:23  */
  assign n5389 = x == 10'b1100000001;
  /* fppowbf16.vhdl:1600:23  */
  assign n5392 = x == 10'b1100000010;
  /* fppowbf16.vhdl:1601:23  */
  assign n5395 = x == 10'b1100000011;
  /* fppowbf16.vhdl:1602:23  */
  assign n5398 = x == 10'b1100000100;
  /* fppowbf16.vhdl:1603:23  */
  assign n5401 = x == 10'b1100000101;
  /* fppowbf16.vhdl:1604:23  */
  assign n5404 = x == 10'b1100000110;
  /* fppowbf16.vhdl:1605:23  */
  assign n5407 = x == 10'b1100000111;
  /* fppowbf16.vhdl:1606:23  */
  assign n5410 = x == 10'b1100001000;
  /* fppowbf16.vhdl:1607:23  */
  assign n5413 = x == 10'b1100001001;
  /* fppowbf16.vhdl:1608:23  */
  assign n5416 = x == 10'b1100001010;
  /* fppowbf16.vhdl:1609:23  */
  assign n5419 = x == 10'b1100001011;
  /* fppowbf16.vhdl:1610:23  */
  assign n5422 = x == 10'b1100001100;
  /* fppowbf16.vhdl:1611:23  */
  assign n5425 = x == 10'b1100001101;
  /* fppowbf16.vhdl:1612:23  */
  assign n5428 = x == 10'b1100001110;
  /* fppowbf16.vhdl:1613:23  */
  assign n5431 = x == 10'b1100001111;
  /* fppowbf16.vhdl:1614:23  */
  assign n5434 = x == 10'b1100010000;
  /* fppowbf16.vhdl:1615:23  */
  assign n5437 = x == 10'b1100010001;
  /* fppowbf16.vhdl:1616:23  */
  assign n5440 = x == 10'b1100010010;
  /* fppowbf16.vhdl:1617:23  */
  assign n5443 = x == 10'b1100010011;
  /* fppowbf16.vhdl:1618:23  */
  assign n5446 = x == 10'b1100010100;
  /* fppowbf16.vhdl:1619:23  */
  assign n5449 = x == 10'b1100010101;
  /* fppowbf16.vhdl:1620:23  */
  assign n5452 = x == 10'b1100010110;
  /* fppowbf16.vhdl:1621:23  */
  assign n5455 = x == 10'b1100010111;
  /* fppowbf16.vhdl:1622:23  */
  assign n5458 = x == 10'b1100011000;
  /* fppowbf16.vhdl:1623:23  */
  assign n5461 = x == 10'b1100011001;
  /* fppowbf16.vhdl:1624:23  */
  assign n5464 = x == 10'b1100011010;
  /* fppowbf16.vhdl:1625:23  */
  assign n5467 = x == 10'b1100011011;
  /* fppowbf16.vhdl:1626:23  */
  assign n5470 = x == 10'b1100011100;
  /* fppowbf16.vhdl:1627:23  */
  assign n5473 = x == 10'b1100011101;
  /* fppowbf16.vhdl:1628:23  */
  assign n5476 = x == 10'b1100011110;
  /* fppowbf16.vhdl:1629:23  */
  assign n5479 = x == 10'b1100011111;
  /* fppowbf16.vhdl:1630:23  */
  assign n5482 = x == 10'b1100100000;
  /* fppowbf16.vhdl:1631:23  */
  assign n5485 = x == 10'b1100100001;
  /* fppowbf16.vhdl:1632:23  */
  assign n5488 = x == 10'b1100100010;
  /* fppowbf16.vhdl:1633:23  */
  assign n5491 = x == 10'b1100100011;
  /* fppowbf16.vhdl:1634:23  */
  assign n5494 = x == 10'b1100100100;
  /* fppowbf16.vhdl:1635:23  */
  assign n5497 = x == 10'b1100100101;
  /* fppowbf16.vhdl:1636:23  */
  assign n5500 = x == 10'b1100100110;
  /* fppowbf16.vhdl:1637:23  */
  assign n5503 = x == 10'b1100100111;
  /* fppowbf16.vhdl:1638:23  */
  assign n5506 = x == 10'b1100101000;
  /* fppowbf16.vhdl:1639:23  */
  assign n5509 = x == 10'b1100101001;
  /* fppowbf16.vhdl:1640:23  */
  assign n5512 = x == 10'b1100101010;
  /* fppowbf16.vhdl:1641:23  */
  assign n5515 = x == 10'b1100101011;
  /* fppowbf16.vhdl:1642:23  */
  assign n5518 = x == 10'b1100101100;
  /* fppowbf16.vhdl:1643:23  */
  assign n5521 = x == 10'b1100101101;
  /* fppowbf16.vhdl:1644:23  */
  assign n5524 = x == 10'b1100101110;
  /* fppowbf16.vhdl:1645:23  */
  assign n5527 = x == 10'b1100101111;
  /* fppowbf16.vhdl:1646:23  */
  assign n5530 = x == 10'b1100110000;
  /* fppowbf16.vhdl:1647:23  */
  assign n5533 = x == 10'b1100110001;
  /* fppowbf16.vhdl:1648:23  */
  assign n5536 = x == 10'b1100110010;
  /* fppowbf16.vhdl:1649:23  */
  assign n5539 = x == 10'b1100110011;
  /* fppowbf16.vhdl:1650:23  */
  assign n5542 = x == 10'b1100110100;
  /* fppowbf16.vhdl:1651:23  */
  assign n5545 = x == 10'b1100110101;
  /* fppowbf16.vhdl:1652:23  */
  assign n5548 = x == 10'b1100110110;
  /* fppowbf16.vhdl:1653:23  */
  assign n5551 = x == 10'b1100110111;
  /* fppowbf16.vhdl:1654:23  */
  assign n5554 = x == 10'b1100111000;
  /* fppowbf16.vhdl:1655:23  */
  assign n5557 = x == 10'b1100111001;
  /* fppowbf16.vhdl:1656:23  */
  assign n5560 = x == 10'b1100111010;
  /* fppowbf16.vhdl:1657:23  */
  assign n5563 = x == 10'b1100111011;
  /* fppowbf16.vhdl:1658:23  */
  assign n5566 = x == 10'b1100111100;
  /* fppowbf16.vhdl:1659:23  */
  assign n5569 = x == 10'b1100111101;
  /* fppowbf16.vhdl:1660:23  */
  assign n5572 = x == 10'b1100111110;
  /* fppowbf16.vhdl:1661:23  */
  assign n5575 = x == 10'b1100111111;
  /* fppowbf16.vhdl:1662:23  */
  assign n5578 = x == 10'b1101000000;
  /* fppowbf16.vhdl:1663:23  */
  assign n5581 = x == 10'b1101000001;
  /* fppowbf16.vhdl:1664:23  */
  assign n5584 = x == 10'b1101000010;
  /* fppowbf16.vhdl:1665:23  */
  assign n5587 = x == 10'b1101000011;
  /* fppowbf16.vhdl:1666:23  */
  assign n5590 = x == 10'b1101000100;
  /* fppowbf16.vhdl:1667:23  */
  assign n5593 = x == 10'b1101000101;
  /* fppowbf16.vhdl:1668:23  */
  assign n5596 = x == 10'b1101000110;
  /* fppowbf16.vhdl:1669:23  */
  assign n5599 = x == 10'b1101000111;
  /* fppowbf16.vhdl:1670:23  */
  assign n5602 = x == 10'b1101001000;
  /* fppowbf16.vhdl:1671:23  */
  assign n5605 = x == 10'b1101001001;
  /* fppowbf16.vhdl:1672:23  */
  assign n5608 = x == 10'b1101001010;
  /* fppowbf16.vhdl:1673:23  */
  assign n5611 = x == 10'b1101001011;
  /* fppowbf16.vhdl:1674:23  */
  assign n5614 = x == 10'b1101001100;
  /* fppowbf16.vhdl:1675:23  */
  assign n5617 = x == 10'b1101001101;
  /* fppowbf16.vhdl:1676:23  */
  assign n5620 = x == 10'b1101001110;
  /* fppowbf16.vhdl:1677:23  */
  assign n5623 = x == 10'b1101001111;
  /* fppowbf16.vhdl:1678:23  */
  assign n5626 = x == 10'b1101010000;
  /* fppowbf16.vhdl:1679:23  */
  assign n5629 = x == 10'b1101010001;
  /* fppowbf16.vhdl:1680:23  */
  assign n5632 = x == 10'b1101010010;
  /* fppowbf16.vhdl:1681:23  */
  assign n5635 = x == 10'b1101010011;
  /* fppowbf16.vhdl:1682:23  */
  assign n5638 = x == 10'b1101010100;
  /* fppowbf16.vhdl:1683:23  */
  assign n5641 = x == 10'b1101010101;
  /* fppowbf16.vhdl:1684:23  */
  assign n5644 = x == 10'b1101010110;
  /* fppowbf16.vhdl:1685:23  */
  assign n5647 = x == 10'b1101010111;
  /* fppowbf16.vhdl:1686:23  */
  assign n5650 = x == 10'b1101011000;
  /* fppowbf16.vhdl:1687:23  */
  assign n5653 = x == 10'b1101011001;
  /* fppowbf16.vhdl:1688:23  */
  assign n5656 = x == 10'b1101011010;
  /* fppowbf16.vhdl:1689:23  */
  assign n5659 = x == 10'b1101011011;
  /* fppowbf16.vhdl:1690:23  */
  assign n5662 = x == 10'b1101011100;
  /* fppowbf16.vhdl:1691:23  */
  assign n5665 = x == 10'b1101011101;
  /* fppowbf16.vhdl:1692:23  */
  assign n5668 = x == 10'b1101011110;
  /* fppowbf16.vhdl:1693:23  */
  assign n5671 = x == 10'b1101011111;
  /* fppowbf16.vhdl:1694:23  */
  assign n5674 = x == 10'b1101100000;
  /* fppowbf16.vhdl:1695:23  */
  assign n5677 = x == 10'b1101100001;
  /* fppowbf16.vhdl:1696:23  */
  assign n5680 = x == 10'b1101100010;
  /* fppowbf16.vhdl:1697:23  */
  assign n5683 = x == 10'b1101100011;
  /* fppowbf16.vhdl:1698:23  */
  assign n5686 = x == 10'b1101100100;
  /* fppowbf16.vhdl:1699:23  */
  assign n5689 = x == 10'b1101100101;
  /* fppowbf16.vhdl:1700:23  */
  assign n5692 = x == 10'b1101100110;
  /* fppowbf16.vhdl:1701:23  */
  assign n5695 = x == 10'b1101100111;
  /* fppowbf16.vhdl:1702:23  */
  assign n5698 = x == 10'b1101101000;
  /* fppowbf16.vhdl:1703:23  */
  assign n5701 = x == 10'b1101101001;
  /* fppowbf16.vhdl:1704:23  */
  assign n5704 = x == 10'b1101101010;
  /* fppowbf16.vhdl:1705:23  */
  assign n5707 = x == 10'b1101101011;
  /* fppowbf16.vhdl:1706:23  */
  assign n5710 = x == 10'b1101101100;
  /* fppowbf16.vhdl:1707:23  */
  assign n5713 = x == 10'b1101101101;
  /* fppowbf16.vhdl:1708:23  */
  assign n5716 = x == 10'b1101101110;
  /* fppowbf16.vhdl:1709:23  */
  assign n5719 = x == 10'b1101101111;
  /* fppowbf16.vhdl:1710:23  */
  assign n5722 = x == 10'b1101110000;
  /* fppowbf16.vhdl:1711:23  */
  assign n5725 = x == 10'b1101110001;
  /* fppowbf16.vhdl:1712:23  */
  assign n5728 = x == 10'b1101110010;
  /* fppowbf16.vhdl:1713:23  */
  assign n5731 = x == 10'b1101110011;
  /* fppowbf16.vhdl:1714:23  */
  assign n5734 = x == 10'b1101110100;
  /* fppowbf16.vhdl:1715:23  */
  assign n5737 = x == 10'b1101110101;
  /* fppowbf16.vhdl:1716:23  */
  assign n5740 = x == 10'b1101110110;
  /* fppowbf16.vhdl:1717:23  */
  assign n5743 = x == 10'b1101110111;
  /* fppowbf16.vhdl:1718:23  */
  assign n5746 = x == 10'b1101111000;
  /* fppowbf16.vhdl:1719:23  */
  assign n5749 = x == 10'b1101111001;
  /* fppowbf16.vhdl:1720:23  */
  assign n5752 = x == 10'b1101111010;
  /* fppowbf16.vhdl:1721:23  */
  assign n5755 = x == 10'b1101111011;
  /* fppowbf16.vhdl:1722:23  */
  assign n5758 = x == 10'b1101111100;
  /* fppowbf16.vhdl:1723:23  */
  assign n5761 = x == 10'b1101111101;
  /* fppowbf16.vhdl:1724:23  */
  assign n5764 = x == 10'b1101111110;
  /* fppowbf16.vhdl:1725:23  */
  assign n5767 = x == 10'b1101111111;
  /* fppowbf16.vhdl:1726:23  */
  assign n5770 = x == 10'b1110000000;
  /* fppowbf16.vhdl:1727:23  */
  assign n5773 = x == 10'b1110000001;
  /* fppowbf16.vhdl:1728:23  */
  assign n5776 = x == 10'b1110000010;
  /* fppowbf16.vhdl:1729:23  */
  assign n5779 = x == 10'b1110000011;
  /* fppowbf16.vhdl:1730:23  */
  assign n5782 = x == 10'b1110000100;
  /* fppowbf16.vhdl:1731:23  */
  assign n5785 = x == 10'b1110000101;
  /* fppowbf16.vhdl:1732:23  */
  assign n5788 = x == 10'b1110000110;
  /* fppowbf16.vhdl:1733:23  */
  assign n5791 = x == 10'b1110000111;
  /* fppowbf16.vhdl:1734:23  */
  assign n5794 = x == 10'b1110001000;
  /* fppowbf16.vhdl:1735:23  */
  assign n5797 = x == 10'b1110001001;
  /* fppowbf16.vhdl:1736:23  */
  assign n5800 = x == 10'b1110001010;
  /* fppowbf16.vhdl:1737:23  */
  assign n5803 = x == 10'b1110001011;
  /* fppowbf16.vhdl:1738:23  */
  assign n5806 = x == 10'b1110001100;
  /* fppowbf16.vhdl:1739:23  */
  assign n5809 = x == 10'b1110001101;
  /* fppowbf16.vhdl:1740:23  */
  assign n5812 = x == 10'b1110001110;
  /* fppowbf16.vhdl:1741:23  */
  assign n5815 = x == 10'b1110001111;
  /* fppowbf16.vhdl:1742:23  */
  assign n5818 = x == 10'b1110010000;
  /* fppowbf16.vhdl:1743:23  */
  assign n5821 = x == 10'b1110010001;
  /* fppowbf16.vhdl:1744:23  */
  assign n5824 = x == 10'b1110010010;
  /* fppowbf16.vhdl:1745:23  */
  assign n5827 = x == 10'b1110010011;
  /* fppowbf16.vhdl:1746:23  */
  assign n5830 = x == 10'b1110010100;
  /* fppowbf16.vhdl:1747:23  */
  assign n5833 = x == 10'b1110010101;
  /* fppowbf16.vhdl:1748:23  */
  assign n5836 = x == 10'b1110010110;
  /* fppowbf16.vhdl:1749:23  */
  assign n5839 = x == 10'b1110010111;
  /* fppowbf16.vhdl:1750:23  */
  assign n5842 = x == 10'b1110011000;
  /* fppowbf16.vhdl:1751:23  */
  assign n5845 = x == 10'b1110011001;
  /* fppowbf16.vhdl:1752:23  */
  assign n5848 = x == 10'b1110011010;
  /* fppowbf16.vhdl:1753:23  */
  assign n5851 = x == 10'b1110011011;
  /* fppowbf16.vhdl:1754:23  */
  assign n5854 = x == 10'b1110011100;
  /* fppowbf16.vhdl:1755:23  */
  assign n5857 = x == 10'b1110011101;
  /* fppowbf16.vhdl:1756:23  */
  assign n5860 = x == 10'b1110011110;
  /* fppowbf16.vhdl:1757:23  */
  assign n5863 = x == 10'b1110011111;
  /* fppowbf16.vhdl:1758:23  */
  assign n5866 = x == 10'b1110100000;
  /* fppowbf16.vhdl:1759:23  */
  assign n5869 = x == 10'b1110100001;
  /* fppowbf16.vhdl:1760:23  */
  assign n5872 = x == 10'b1110100010;
  /* fppowbf16.vhdl:1761:23  */
  assign n5875 = x == 10'b1110100011;
  /* fppowbf16.vhdl:1762:23  */
  assign n5878 = x == 10'b1110100100;
  /* fppowbf16.vhdl:1763:23  */
  assign n5881 = x == 10'b1110100101;
  /* fppowbf16.vhdl:1764:23  */
  assign n5884 = x == 10'b1110100110;
  /* fppowbf16.vhdl:1765:23  */
  assign n5887 = x == 10'b1110100111;
  /* fppowbf16.vhdl:1766:23  */
  assign n5890 = x == 10'b1110101000;
  /* fppowbf16.vhdl:1767:23  */
  assign n5893 = x == 10'b1110101001;
  /* fppowbf16.vhdl:1768:23  */
  assign n5896 = x == 10'b1110101010;
  /* fppowbf16.vhdl:1769:23  */
  assign n5899 = x == 10'b1110101011;
  /* fppowbf16.vhdl:1770:23  */
  assign n5902 = x == 10'b1110101100;
  /* fppowbf16.vhdl:1771:23  */
  assign n5905 = x == 10'b1110101101;
  /* fppowbf16.vhdl:1772:23  */
  assign n5908 = x == 10'b1110101110;
  /* fppowbf16.vhdl:1773:23  */
  assign n5911 = x == 10'b1110101111;
  /* fppowbf16.vhdl:1774:23  */
  assign n5914 = x == 10'b1110110000;
  /* fppowbf16.vhdl:1775:23  */
  assign n5917 = x == 10'b1110110001;
  /* fppowbf16.vhdl:1776:23  */
  assign n5920 = x == 10'b1110110010;
  /* fppowbf16.vhdl:1777:23  */
  assign n5923 = x == 10'b1110110011;
  /* fppowbf16.vhdl:1778:23  */
  assign n5926 = x == 10'b1110110100;
  /* fppowbf16.vhdl:1779:23  */
  assign n5929 = x == 10'b1110110101;
  /* fppowbf16.vhdl:1780:23  */
  assign n5932 = x == 10'b1110110110;
  /* fppowbf16.vhdl:1781:23  */
  assign n5935 = x == 10'b1110110111;
  /* fppowbf16.vhdl:1782:23  */
  assign n5938 = x == 10'b1110111000;
  /* fppowbf16.vhdl:1783:23  */
  assign n5941 = x == 10'b1110111001;
  /* fppowbf16.vhdl:1784:23  */
  assign n5944 = x == 10'b1110111010;
  /* fppowbf16.vhdl:1785:23  */
  assign n5947 = x == 10'b1110111011;
  /* fppowbf16.vhdl:1786:23  */
  assign n5950 = x == 10'b1110111100;
  /* fppowbf16.vhdl:1787:23  */
  assign n5953 = x == 10'b1110111101;
  /* fppowbf16.vhdl:1788:23  */
  assign n5956 = x == 10'b1110111110;
  /* fppowbf16.vhdl:1789:23  */
  assign n5959 = x == 10'b1110111111;
  /* fppowbf16.vhdl:1790:23  */
  assign n5962 = x == 10'b1111000000;
  /* fppowbf16.vhdl:1791:23  */
  assign n5965 = x == 10'b1111000001;
  /* fppowbf16.vhdl:1792:23  */
  assign n5968 = x == 10'b1111000010;
  /* fppowbf16.vhdl:1793:23  */
  assign n5971 = x == 10'b1111000011;
  /* fppowbf16.vhdl:1794:23  */
  assign n5974 = x == 10'b1111000100;
  /* fppowbf16.vhdl:1795:23  */
  assign n5977 = x == 10'b1111000101;
  /* fppowbf16.vhdl:1796:23  */
  assign n5980 = x == 10'b1111000110;
  /* fppowbf16.vhdl:1797:23  */
  assign n5983 = x == 10'b1111000111;
  /* fppowbf16.vhdl:1798:23  */
  assign n5986 = x == 10'b1111001000;
  /* fppowbf16.vhdl:1799:23  */
  assign n5989 = x == 10'b1111001001;
  /* fppowbf16.vhdl:1800:23  */
  assign n5992 = x == 10'b1111001010;
  /* fppowbf16.vhdl:1801:23  */
  assign n5995 = x == 10'b1111001011;
  /* fppowbf16.vhdl:1802:23  */
  assign n5998 = x == 10'b1111001100;
  /* fppowbf16.vhdl:1803:23  */
  assign n6001 = x == 10'b1111001101;
  /* fppowbf16.vhdl:1804:23  */
  assign n6004 = x == 10'b1111001110;
  /* fppowbf16.vhdl:1805:23  */
  assign n6007 = x == 10'b1111001111;
  /* fppowbf16.vhdl:1806:23  */
  assign n6010 = x == 10'b1111010000;
  /* fppowbf16.vhdl:1807:23  */
  assign n6013 = x == 10'b1111010001;
  /* fppowbf16.vhdl:1808:23  */
  assign n6016 = x == 10'b1111010010;
  /* fppowbf16.vhdl:1809:23  */
  assign n6019 = x == 10'b1111010011;
  /* fppowbf16.vhdl:1810:23  */
  assign n6022 = x == 10'b1111010100;
  /* fppowbf16.vhdl:1811:23  */
  assign n6025 = x == 10'b1111010101;
  /* fppowbf16.vhdl:1812:23  */
  assign n6028 = x == 10'b1111010110;
  /* fppowbf16.vhdl:1813:23  */
  assign n6031 = x == 10'b1111010111;
  /* fppowbf16.vhdl:1814:23  */
  assign n6034 = x == 10'b1111011000;
  /* fppowbf16.vhdl:1815:23  */
  assign n6037 = x == 10'b1111011001;
  /* fppowbf16.vhdl:1816:23  */
  assign n6040 = x == 10'b1111011010;
  /* fppowbf16.vhdl:1817:23  */
  assign n6043 = x == 10'b1111011011;
  /* fppowbf16.vhdl:1818:23  */
  assign n6046 = x == 10'b1111011100;
  /* fppowbf16.vhdl:1819:23  */
  assign n6049 = x == 10'b1111011101;
  /* fppowbf16.vhdl:1820:23  */
  assign n6052 = x == 10'b1111011110;
  /* fppowbf16.vhdl:1821:23  */
  assign n6055 = x == 10'b1111011111;
  /* fppowbf16.vhdl:1822:23  */
  assign n6058 = x == 10'b1111100000;
  /* fppowbf16.vhdl:1823:23  */
  assign n6061 = x == 10'b1111100001;
  /* fppowbf16.vhdl:1824:23  */
  assign n6064 = x == 10'b1111100010;
  /* fppowbf16.vhdl:1825:23  */
  assign n6067 = x == 10'b1111100011;
  /* fppowbf16.vhdl:1826:23  */
  assign n6070 = x == 10'b1111100100;
  /* fppowbf16.vhdl:1827:23  */
  assign n6073 = x == 10'b1111100101;
  /* fppowbf16.vhdl:1828:23  */
  assign n6076 = x == 10'b1111100110;
  /* fppowbf16.vhdl:1829:23  */
  assign n6079 = x == 10'b1111100111;
  /* fppowbf16.vhdl:1830:23  */
  assign n6082 = x == 10'b1111101000;
  /* fppowbf16.vhdl:1831:23  */
  assign n6085 = x == 10'b1111101001;
  /* fppowbf16.vhdl:1832:23  */
  assign n6088 = x == 10'b1111101010;
  /* fppowbf16.vhdl:1833:23  */
  assign n6091 = x == 10'b1111101011;
  /* fppowbf16.vhdl:1834:23  */
  assign n6094 = x == 10'b1111101100;
  /* fppowbf16.vhdl:1835:23  */
  assign n6097 = x == 10'b1111101101;
  /* fppowbf16.vhdl:1836:23  */
  assign n6100 = x == 10'b1111101110;
  /* fppowbf16.vhdl:1837:23  */
  assign n6103 = x == 10'b1111101111;
  /* fppowbf16.vhdl:1838:23  */
  assign n6106 = x == 10'b1111110000;
  /* fppowbf16.vhdl:1839:23  */
  assign n6109 = x == 10'b1111110001;
  /* fppowbf16.vhdl:1840:23  */
  assign n6112 = x == 10'b1111110010;
  /* fppowbf16.vhdl:1841:23  */
  assign n6115 = x == 10'b1111110011;
  /* fppowbf16.vhdl:1842:23  */
  assign n6118 = x == 10'b1111110100;
  /* fppowbf16.vhdl:1843:23  */
  assign n6121 = x == 10'b1111110101;
  /* fppowbf16.vhdl:1844:23  */
  assign n6124 = x == 10'b1111110110;
  /* fppowbf16.vhdl:1845:23  */
  assign n6127 = x == 10'b1111110111;
  /* fppowbf16.vhdl:1846:23  */
  assign n6130 = x == 10'b1111111000;
  /* fppowbf16.vhdl:1847:23  */
  assign n6133 = x == 10'b1111111001;
  /* fppowbf16.vhdl:1848:23  */
  assign n6136 = x == 10'b1111111010;
  /* fppowbf16.vhdl:1849:23  */
  assign n6139 = x == 10'b1111111011;
  /* fppowbf16.vhdl:1850:23  */
  assign n6142 = x == 10'b1111111100;
  /* fppowbf16.vhdl:1851:23  */
  assign n6145 = x == 10'b1111111101;
  /* fppowbf16.vhdl:1852:23  */
  assign n6148 = x == 10'b1111111110;
  /* fppowbf16.vhdl:1853:23  */
  assign n6151 = x == 10'b1111111111;
  assign n6153 = {n6151, n6148, n6145, n6142, n6139, n6136, n6133, n6130, n6127, n6124, n6121, n6118, n6115, n6112, n6109, n6106, n6103, n6100, n6097, n6094, n6091, n6088, n6085, n6082, n6079, n6076, n6073, n6070, n6067, n6064, n6061, n6058, n6055, n6052, n6049, n6046, n6043, n6040, n6037, n6034, n6031, n6028, n6025, n6022, n6019, n6016, n6013, n6010, n6007, n6004, n6001, n5998, n5995, n5992, n5989, n5986, n5983, n5980, n5977, n5974, n5971, n5968, n5965, n5962, n5959, n5956, n5953, n5950, n5947, n5944, n5941, n5938, n5935, n5932, n5929, n5926, n5923, n5920, n5917, n5914, n5911, n5908, n5905, n5902, n5899, n5896, n5893, n5890, n5887, n5884, n5881, n5878, n5875, n5872, n5869, n5866, n5863, n5860, n5857, n5854, n5851, n5848, n5845, n5842, n5839, n5836, n5833, n5830, n5827, n5824, n5821, n5818, n5815, n5812, n5809, n5806, n5803, n5800, n5797, n5794, n5791, n5788, n5785, n5782, n5779, n5776, n5773, n5770, n5767, n5764, n5761, n5758, n5755, n5752, n5749, n5746, n5743, n5740, n5737, n5734, n5731, n5728, n5725, n5722, n5719, n5716, n5713, n5710, n5707, n5704, n5701, n5698, n5695, n5692, n5689, n5686, n5683, n5680, n5677, n5674, n5671, n5668, n5665, n5662, n5659, n5656, n5653, n5650, n5647, n5644, n5641, n5638, n5635, n5632, n5629, n5626, n5623, n5620, n5617, n5614, n5611, n5608, n5605, n5602, n5599, n5596, n5593, n5590, n5587, n5584, n5581, n5578, n5575, n5572, n5569, n5566, n5563, n5560, n5557, n5554, n5551, n5548, n5545, n5542, n5539, n5536, n5533, n5530, n5527, n5524, n5521, n5518, n5515, n5512, n5509, n5506, n5503, n5500, n5497, n5494, n5491, n5488, n5485, n5482, n5479, n5476, n5473, n5470, n5467, n5464, n5461, n5458, n5455, n5452, n5449, n5446, n5443, n5440, n5437, n5434, n5431, n5428, n5425, n5422, n5419, n5416, n5413, n5410, n5407, n5404, n5401, n5398, n5395, n5392, n5389, n5386, n5383, n5380, n5377, n5374, n5371, n5368, n5365, n5362, n5359, n5356, n5353, n5350, n5347, n5344, n5341, n5338, n5335, n5332, n5329, n5326, n5323, n5320, n5317, n5314, n5311, n5308, n5305, n5302, n5299, n5296, n5293, n5290, n5287, n5284, n5281, n5278, n5275, n5272, n5269, n5266, n5263, n5260, n5257, n5254, n5251, n5248, n5245, n5242, n5239, n5236, n5233, n5230, n5227, n5224, n5221, n5218, n5215, n5212, n5209, n5206, n5203, n5200, n5197, n5194, n5191, n5188, n5185, n5182, n5179, n5176, n5173, n5170, n5167, n5164, n5161, n5158, n5155, n5152, n5149, n5146, n5143, n5140, n5137, n5134, n5131, n5128, n5125, n5122, n5119, n5116, n5113, n5110, n5107, n5104, n5101, n5098, n5095, n5092, n5089, n5086, n5083, n5080, n5077, n5074, n5071, n5068, n5065, n5062, n5059, n5056, n5053, n5050, n5047, n5044, n5041, n5038, n5035, n5032, n5029, n5026, n5023, n5020, n5017, n5014, n5011, n5008, n5005, n5002, n4999, n4996, n4993, n4990, n4987, n4984, n4981, n4978, n4975, n4972, n4969, n4966, n4963, n4960, n4957, n4954, n4951, n4948, n4945, n4942, n4939, n4936, n4933, n4930, n4927, n4924, n4921, n4918, n4915, n4912, n4909, n4906, n4903, n4900, n4897, n4894, n4891, n4888, n4885, n4882, n4879, n4876, n4873, n4870, n4867, n4864, n4861, n4858, n4855, n4852, n4849, n4846, n4843, n4840, n4837, n4834, n4831, n4828, n4825, n4822, n4819, n4816, n4813, n4810, n4807, n4804, n4801, n4798, n4795, n4792, n4789, n4786, n4783, n4780, n4777, n4774, n4771, n4768, n4765, n4762, n4759, n4756, n4753, n4750, n4747, n4744, n4741, n4738, n4735, n4732, n4729, n4726, n4723, n4720, n4717, n4714, n4711, n4708, n4705, n4702, n4699, n4696, n4693, n4690, n4687, n4684, n4681, n4678, n4675, n4672, n4669, n4666, n4663, n4660, n4657, n4654, n4651, n4648, n4645, n4642, n4639, n4636, n4633, n4630, n4627, n4624, n4621, n4618, n4615, n4612, n4609, n4606, n4603, n4600, n4597, n4594, n4591, n4588, n4585, n4582, n4579, n4576, n4573, n4570, n4567, n4564, n4561, n4558, n4555, n4552, n4549, n4546, n4543, n4540, n4537, n4534, n4531, n4528, n4525, n4522, n4519, n4516, n4513, n4510, n4507, n4504, n4501, n4498, n4495, n4492, n4489, n4486, n4483, n4480, n4477, n4474, n4471, n4468, n4465, n4462, n4459, n4456, n4453, n4450, n4447, n4444, n4441, n4438, n4435, n4432, n4429, n4426, n4423, n4420, n4417, n4414, n4411, n4408, n4405, n4402, n4399, n4396, n4393, n4390, n4387, n4384, n4381, n4378, n4375, n4372, n4369, n4366, n4363, n4360, n4357, n4354, n4351, n4348, n4345, n4342, n4339, n4336, n4333, n4330, n4327, n4324, n4321, n4318, n4315, n4312, n4309, n4306, n4303, n4300, n4297, n4294, n4291, n4288, n4285, n4282, n4279, n4276, n4273, n4270, n4267, n4264, n4261, n4258, n4255, n4252, n4249, n4246, n4243, n4240, n4237, n4234, n4231, n4228, n4225, n4222, n4219, n4216, n4213, n4210, n4207, n4204, n4201, n4198, n4195, n4192, n4189, n4186, n4183, n4180, n4177, n4174, n4171, n4168, n4165, n4162, n4159, n4156, n4153, n4150, n4147, n4144, n4141, n4138, n4135, n4132, n4129, n4126, n4123, n4120, n4117, n4114, n4111, n4108, n4105, n4102, n4099, n4096, n4093, n4090, n4087, n4084, n4081, n4078, n4075, n4072, n4069, n4066, n4063, n4060, n4057, n4054, n4051, n4048, n4045, n4042, n4039, n4036, n4033, n4030, n4027, n4024, n4021, n4018, n4015, n4012, n4009, n4006, n4003, n4000, n3997, n3994, n3991, n3988, n3985, n3982, n3979, n3976, n3973, n3970, n3967, n3964, n3961, n3958, n3955, n3952, n3949, n3946, n3943, n3940, n3937, n3934, n3931, n3928, n3925, n3922, n3919, n3916, n3913, n3910, n3907, n3904, n3901, n3898, n3895, n3892, n3889, n3886, n3883, n3880, n3877, n3874, n3871, n3868, n3865, n3862, n3859, n3856, n3853, n3850, n3847, n3844, n3841, n3838, n3835, n3832, n3829, n3826, n3823, n3820, n3817, n3814, n3811, n3808, n3805, n3802, n3799, n3796, n3793, n3790, n3787, n3784, n3781, n3778, n3775, n3772, n3769, n3766, n3763, n3760, n3757, n3754, n3751, n3748, n3745, n3742, n3739, n3736, n3733, n3730, n3727, n3724, n3721, n3718, n3715, n3712, n3709, n3706, n3703, n3700, n3697, n3694, n3691, n3688, n3685, n3682, n3679, n3676, n3673, n3670, n3667, n3664, n3661, n3658, n3655, n3652, n3649, n3646, n3643, n3640, n3637, n3634, n3631, n3628, n3625, n3622, n3619, n3616, n3613, n3610, n3607, n3604, n3601, n3598, n3595, n3592, n3589, n3586, n3583, n3580, n3577, n3574, n3571, n3568, n3565, n3562, n3559, n3556, n3553, n3550, n3547, n3544, n3541, n3538, n3535, n3532, n3529, n3526, n3523, n3520, n3517, n3514, n3511, n3508, n3505, n3502, n3499, n3496, n3493, n3490, n3487, n3484, n3481, n3478, n3475, n3472, n3469, n3466, n3463, n3460, n3457, n3454, n3451, n3448, n3445, n3442, n3439, n3436, n3433, n3430, n3427, n3424, n3421, n3418, n3415, n3412, n3409, n3406, n3403, n3400, n3397, n3394, n3391, n3388, n3385, n3382, n3379, n3376, n3373, n3370, n3367, n3364, n3361, n3358, n3355, n3352, n3349, n3346, n3343, n3340, n3337, n3334, n3331, n3328, n3325, n3322, n3319, n3316, n3313, n3310, n3307, n3304, n3301, n3298, n3295, n3292, n3289, n3286, n3283, n3280, n3277, n3274, n3271, n3268, n3265, n3262, n3259, n3256, n3253, n3250, n3247, n3244, n3241, n3238, n3235, n3232, n3229, n3226, n3223, n3220, n3217, n3214, n3211, n3208, n3205, n3202, n3199, n3196, n3193, n3190, n3187, n3184, n3181, n3178, n3175, n3172, n3169, n3166, n3163, n3160, n3157, n3154, n3151, n3148, n3145, n3142, n3139, n3136, n3133, n3130, n3127, n3124, n3121, n3118, n3115, n3112, n3109, n3106, n3103, n3100, n3097, n3094, n3091, n3088, n3085, n3082};
  /* fppowbf16.vhdl:829:4  */
  always @*
    case (n6153)
      1024'b1000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0111111111100;
      1024'b0100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0111111111000;
      1024'b0010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0111111110100;
      1024'b0001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0111111110000;
      1024'b0000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0111111101100;
      1024'b0000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0111111101000;
      1024'b0000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0111111100100;
      1024'b0000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0111111100000;
      1024'b0000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0111111011100;
      1024'b0000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0111111011000;
      1024'b0000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0111111010100;
      1024'b0000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0111111010000;
      1024'b0000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0111111001100;
      1024'b0000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0111111001000;
      1024'b0000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0111111000100;
      1024'b0000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0111111000000;
      1024'b0000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0111110111101;
      1024'b0000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0111110111001;
      1024'b0000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0111110110101;
      1024'b0000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0111110110001;
      1024'b0000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0111110101101;
      1024'b0000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0111110101001;
      1024'b0000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0111110100101;
      1024'b0000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0111110100001;
      1024'b0000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0111110011101;
      1024'b0000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0111110011001;
      1024'b0000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0111110010101;
      1024'b0000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0111110010010;
      1024'b0000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0111110001110;
      1024'b0000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0111110001010;
      1024'b0000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0111110000110;
      1024'b0000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0111110000010;
      1024'b0000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0111101111110;
      1024'b0000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0111101111010;
      1024'b0000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0111101110110;
      1024'b0000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0111101110011;
      1024'b0000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0111101101111;
      1024'b0000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0111101101011;
      1024'b0000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0111101100111;
      1024'b0000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0111101100011;
      1024'b0000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0111101011111;
      1024'b0000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0111101011011;
      1024'b0000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0111101011000;
      1024'b0000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0111101010100;
      1024'b0000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0111101010000;
      1024'b0000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0111101001100;
      1024'b0000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0111101001000;
      1024'b0000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0111101000100;
      1024'b0000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0111101000001;
      1024'b0000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0111100111101;
      1024'b0000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0111100111001;
      1024'b0000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0111100110101;
      1024'b0000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0111100110001;
      1024'b0000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0111100101110;
      1024'b0000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0111100101010;
      1024'b0000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0111100100110;
      1024'b0000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0111100100010;
      1024'b0000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0111100011110;
      1024'b0000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0111100011011;
      1024'b0000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0111100010111;
      1024'b0000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0111100010011;
      1024'b0000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0111100001111;
      1024'b0000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0111100001100;
      1024'b0000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0111100001000;
      1024'b0000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0111100000100;
      1024'b0000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0111100000000;
      1024'b0000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0111011111101;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0111011111001;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0111011110101;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0111011110001;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0111011101110;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0111011101010;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0111011100110;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0111011100010;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0111011011111;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0111011011011;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0111011010111;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0111011010100;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0111011010000;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0111011001100;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0111011001000;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0111011000101;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0111011000001;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0111010111101;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0111010111010;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0111010110110;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0111010110010;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0111010101111;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0111010101011;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0111010100111;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0111010100100;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0111010100000;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0111010011100;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0111010011001;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0111010010101;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0111010010001;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0111010001110;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0111010001010;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0111010000111;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0111010000011;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0111001111111;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0111001111100;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0111001111000;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0111001110100;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0111001110001;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0111001101101;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0111001101010;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0111001100110;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0111001100010;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0111001011111;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0111001011011;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0111001011000;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0111001010100;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0111001010000;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0111001001101;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0111001001001;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0111001000110;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0111001000010;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0111000111111;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0111000111011;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0111000111000;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0111000110100;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0111000110000;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0111000101101;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0111000101001;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0111000100110;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0111000100010;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0111000011111;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0111000011011;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0111000011000;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0111000010100;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0111000010001;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0111000001101;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0111000001010;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0111000000110;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0111000000011;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0110111111111;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0110111111100;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0110111111000;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0110111110101;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0110111110001;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0110111101110;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0110111101010;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0110111100111;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0110111100011;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0110111100000;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0110111011100;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0110111011001;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0110111010101;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0110111010010;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0110111001110;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0110111001011;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0110111001000;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0110111000100;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0110111000001;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0110110111101;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0110110111010;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0110110110110;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0110110110011;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0110110101111;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0110110101100;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0110110101001;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0110110100101;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0110110100010;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0110110011110;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0110110011011;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0110110011000;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0110110010100;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0110110010001;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0110110001101;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0110110001010;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0110110000111;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0110110000011;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0110110000000;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0110101111101;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0110101111001;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0110101110110;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0110101110010;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0110101101111;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0110101101100;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0110101101000;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0110101100101;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0110101100010;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0110101011110;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0110101011011;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0110101011000;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0110101010100;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0110101010001;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0110101001110;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0110101001010;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0110101000111;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0110101000100;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0110101000000;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0110100111101;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0110100111010;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0110100110110;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0110100110011;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0110100110000;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0110100101101;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0110100101001;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0110100100110;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0110100100011;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0110100011111;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0110100011100;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0110100011001;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0110100010110;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0110100010010;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0110100001111;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0110100001100;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0110100001001;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0110100000101;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0110100000010;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0110011111111;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0110011111100;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0110011111000;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0110011110101;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0110011110010;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0110011101111;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0110011101011;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0110011101000;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0110011100101;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0110011100010;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0110011011110;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0110011011011;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0110011011000;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0110011010101;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0110011010010;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0110011001110;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0110011001011;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0110011001000;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0110011000101;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0110011000010;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0110010111110;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0110010111011;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0110010111000;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0110010110101;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0110010110010;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0110010101111;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0110010101011;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0110010101000;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0110010100101;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0110010100010;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0110010011111;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0110010011100;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0110010011000;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0110010010101;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0110010010010;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0110010001111;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0110010001100;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0110010001001;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0110010000110;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0110010000010;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0110001111111;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0110001111100;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0110001111001;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0110001110110;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0110001110011;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0110001110000;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0110001101101;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0110001101010;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0110001100110;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0110001100011;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0110001100000;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0110001011101;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0110001011010;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0110001010111;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0110001010100;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0110001010001;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0110001001110;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0110001001011;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0110001001000;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0110001000101;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0110001000001;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0110000111110;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0110000111011;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0110000111000;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0110000110101;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0110000110010;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0110000101111;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0110000101100;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0110000101001;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0110000100110;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0110000100011;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0110000100000;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0110000011101;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0110000011010;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0110000010111;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0110000010100;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0110000010001;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0110000001110;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0110000001011;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0110000001000;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0110000000101;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0110000000010;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0101111111111;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0101111111100;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0101111111001;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0101111110110;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0101111110011;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0101111110000;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0101111101101;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0101111101010;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0101111100111;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0101111100100;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0101111100001;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0101111011110;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0101111011011;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0101111011000;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0101111010101;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0101111010010;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0101111001111;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0101111001100;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0101111001001;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0101111000110;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0101111000011;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0101111000000;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0101110111101;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0101110111011;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0101110111000;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0101110110101;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0101110110010;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0101110101111;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0101110101100;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0101110101001;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0101110100110;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0101110100011;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0101110100000;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0101110011101;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0101110011010;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0101110011000;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0101110010101;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0101110010010;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0101110001111;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0101110001100;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0101110001001;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0101110000110;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0101110000011;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0101110000000;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0101101111110;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0101101111011;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0101101111000;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0101101110101;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0101101110010;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0101101101111;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0101101101100;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0101101101010;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0101101100111;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0101101100100;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0101101100001;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0101101011110;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0101101011011;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0101101011000;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0101101010110;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0101101010011;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0101101010000;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0101101001101;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0101101001010;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0101101001000;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0101101000101;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0101101000010;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0101100111111;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0101100111100;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0101100111001;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0101100110111;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0101100110100;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0101100110001;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0101100101110;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0101100101011;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0101100101001;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0101100100110;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0101100100011;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0101100100000;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0101100011110;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0101100011011;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0101100011000;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0101100010101;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0101100010010;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0101100010000;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0101100001101;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0101100001010;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0101100000111;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0101100000101;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0101100000010;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0101011111111;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0101011111100;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0101011111010;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0101011110111;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0101011110100;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0101011110001;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0101011101111;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0101011101100;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0101011101001;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0101011100111;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0101011100100;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0101011100001;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0101011011110;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0101011011100;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0101011011001;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0101011010110;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0101011010011;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0101011010001;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0101011001110;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0101011001011;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0101011001001;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0101011000110;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0101011000011;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0101011000001;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0101010111110;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0101010111011;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0101010111001;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0101010110110;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0101010110011;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0101010110001;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0101010101110;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0101010101011;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0101010101001;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0101010100110;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0101010100011;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0101010100001;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0101010011110;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0101010011011;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0101010011001;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0101010010110;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0101010010011;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0101010010001;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0101010001110;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0101010001011;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0101010001001;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0101010000110;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0101010000011;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0101010000001;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0101001111110;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0101001111100;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0101001111001;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0101001110110;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0101001110100;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0101001110001;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0101001101111;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0101001101100;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0101001101001;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0101001100111;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0101001100100;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0101001100010;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0101001011111;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0101001011100;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0101001011010;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0101001010111;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0101001010101;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0101001010010;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0101001001111;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0101001001101;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0101001001010;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0101001001000;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0101001000101;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0101001000011;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0101001000000;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0101000111101;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0101000111011;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0101000111000;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0101000110110;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0101000110011;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0101000110001;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0101000101110;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0101000101100;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0101000101001;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0101000100110;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0101000100100;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0101000100001;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0101000011111;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0101000011100;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0101000011010;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0101000010111;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0101000010101;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0101000010010;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0101000010000;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0101000001101;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0101000001011;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0101000001000;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0101000000110;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0101000000011;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0101000000001;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0100111111110;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0100111111100;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0100111111001;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0100111110111;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0100111110100;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0100111110010;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0100111101111;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0100111101101;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0100111101010;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0100111101000;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0100111100101;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0100111100011;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0100111100000;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0100111011110;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0100111011011;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0100111011001;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0100111010111;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0100111010100;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0100111010010;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0100111001111;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0100111001101;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0100111001010;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0100111001000;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0100111000101;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0100111000011;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0100111000001;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0100110111110;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0100110111100;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0100110111001;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0100110110111;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b0100110110100;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1101001011011;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1101001010100;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1101001001101;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1101001000111;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1101001000000;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1101000111010;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1101000110011;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1101000101101;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1101000100110;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1101000100000;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1101000011001;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1101000010010;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1101000001100;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1101000000101;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1100111111111;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1100111111000;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1100111110010;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1100111101011;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1100111100101;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1100111011111;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1100111011000;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1100111010010;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1100111001011;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1100111000101;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1100110111110;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1100110111000;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1100110110001;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1100110101011;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1100110100101;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1100110011110;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1100110011000;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1100110010001;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1100110001011;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1100110000101;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1100101111110;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1100101111000;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1100101110010;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1100101101011;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1100101100101;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1100101011110;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1100101011000;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1100101010010;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1100101001011;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1100101000101;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1100100111111;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1100100111001;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1100100110010;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1100100101100;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1100100100110;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1100100011111;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1100100011001;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1100100010011;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1100100001101;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1100100000110;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1100100000000;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1100011111010;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1100011110100;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1100011101101;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1100011100111;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1100011100001;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1100011011011;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1100011010100;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1100011001110;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1100011001000;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1100011000010;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1100010111100;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1100010110101;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1100010101111;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1100010101001;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1100010100011;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1100010011101;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1100010010111;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1100010010000;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1100010001010;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1100010000100;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1100001111110;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1100001111000;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1100001110010;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1100001101100;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1100001100110;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1100001100000;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1100001011001;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1100001010011;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1100001001101;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1100001000111;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1100001000001;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1100000111011;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1100000110101;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1100000101111;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1100000101001;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1100000100011;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1100000011101;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1100000010111;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1100000010001;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1100000001011;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1100000000101;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1011111111111;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1011111111001;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1011111110011;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1011111101101;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1011111100111;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1011111100001;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1011111011011;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1011111010101;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1011111001111;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1011111001001;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1011111000011;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1011110111101;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1011110110111;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1011110110001;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1011110101011;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1011110100101;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1011110100000;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1011110011010;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1011110010100;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1011110001110;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1011110001000;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1011110000010;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1011101111100;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1011101110110;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1011101110001;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1011101101011;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1011101100101;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1011101011111;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1011101011001;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1011101010011;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1011101001101;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1011101001000;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1011101000010;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1011100111100;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1011100110110;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1011100110000;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1011100101011;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1011100100101;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1011100011111;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1011100011001;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1011100010011;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1011100001110;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1011100001000;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1011100000010;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1011011111100;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1011011110111;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1011011110001;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1011011101011;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1011011100110;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1011011100000;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1011011011010;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1011011010100;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1011011001111;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1011011001001;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1011011000011;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1011010111110;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1011010111000;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1011010110010;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1011010101101;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1011010100111;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1011010100001;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1011010011100;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1011010010110;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1011010010000;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1011010001011;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1011010000101;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1011001111111;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1011001111010;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1011001110100;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1011001101111;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1011001101001;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1011001100011;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1011001011110;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1011001011000;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1011001010011;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1011001001101;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1011001000111;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1011001000010;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1011000111100;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1011000110111;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1011000110001;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1011000101100;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1011000100110;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1011000100001;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1011000011011;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1011000010110;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1011000010000;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1011000001010;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1011000000101;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1010111111111;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1010111111010;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1010111110100;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1010111101111;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1010111101010;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1010111100100;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1010111011111;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1010111011001;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1010111010100;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1010111001110;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1010111001001;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1010111000011;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1010110111110;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1010110111000;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1010110110011;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1010110101110;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1010110101000;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1010110100011;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1010110011101;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1010110011000;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1010110010011;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1010110001101;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1010110001000;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1010110000010;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1010101111101;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1010101111000;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1010101110010;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1010101101101;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1010101101000;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1010101100010;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1010101011101;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1010101011000;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1010101010010;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1010101001101;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1010101001000;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1010101000010;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1010100111101;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1010100111000;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1010100110010;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1010100101101;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1010100101000;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1010100100010;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1010100011101;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1010100011000;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1010100010011;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1010100001101;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1010100001000;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1010100000011;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1010011111110;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1010011111000;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1010011110011;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1010011101110;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1010011101001;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1010011100011;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1010011011110;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1010011011001;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1010011010100;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1010011001111;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1010011001001;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1010011000100;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1010010111111;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1010010111010;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1010010110101;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1010010101111;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1010010101010;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1010010100101;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1010010100000;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1010010011011;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1010010010110;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1010010010001;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1010010001011;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1010010000110;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1010010000001;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1010001111100;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1010001110111;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1010001110010;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1010001101101;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1010001101000;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1010001100010;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1010001011101;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1010001011000;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1010001010011;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1010001001110;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1010001001001;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1010001000100;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1010000111111;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1010000111010;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1010000110101;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1010000110000;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1010000101011;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1010000100110;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1010000100001;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1010000011100;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1010000010111;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1010000010010;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1010000001101;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1010000001000;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1010000000011;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1001111111110;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1001111111001;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1001111110100;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1001111101111;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1001111101010;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1001111100101;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1001111100000;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1001111011011;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1001111010110;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1001111010001;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1001111001100;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1001111000111;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1001111000010;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1001110111101;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1001110111000;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1001110110011;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1001110101110;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1001110101001;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1001110100100;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1001110011111;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1001110011011;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1001110010110;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1001110010001;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1001110001100;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1001110000111;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1001110000010;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1001101111101;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1001101111000;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1001101110011;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1001101101111;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1001101101010;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1001101100101;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1001101100000;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1001101011011;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1001101010110;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1001101010010;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1001101001101;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1001101001000;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1001101000011;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1001100111110;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1001100111001;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1001100110101;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1001100110000;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1001100101011;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1001100100110;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1001100100001;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1001100011101;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1001100011000;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1001100010011;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1001100001110;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1001100001010;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1001100000101;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1001100000000;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1001011111011;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1001011110111;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1001011110010;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1001011101101;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1001011101000;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1001011100100;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1001011011111;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1001011011010;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1001011010110;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1001011010001;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1001011001100;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1001011000111;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1001011000011;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1001010111110;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1001010111001;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1001010110101;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1001010110000;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1001010101011;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1001010100111;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1001010100010;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1001010011101;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1001010011001;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1001010010100;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1001010001111;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1001010001011;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1001010000110;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1001010000010;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1001001111101;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1001001111000;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1001001110100;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1001001101111;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1001001101010;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1001001100110;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1001001100001;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1001001011101;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1001001011000;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1001001010100;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1001001001111;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1001001001010;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1001001000110;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1001001000001;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1001000111101;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1001000111000;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1001000110100;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1001000101111;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1001000101010;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1001000100110;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1001000100001;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1001000011101;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1001000011000;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1001000010100;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1001000001111;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1001000001011;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1001000000110;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1001000000010;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1000111111101;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1000111111001;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1000111110100;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1000111110000;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1000111101011;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1000111100111;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1000111100010;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1000111011110;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1000111011001;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1000111010101;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1000111010001;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1000111001100;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1000111001000;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1000111000011;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1000110111111;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1000110111010;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1000110110110;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1000110110001;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1000110101101;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1000110101001;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1000110100100;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1000110100000;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1000110011011;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1000110010111;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1000110010011;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1000110001110;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1000110001010;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1000110000101;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1000110000001;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1000101111101;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1000101111000;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1000101110100;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1000101110000;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1000101101011;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1000101100111;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1000101100011;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1000101011110;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1000101011010;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1000101010101;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1000101010001;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1000101001101;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1000101001001;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1000101000100;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1000101000000;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1000100111100;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1000100110111;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1000100110011;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1000100101111;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1000100101010;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1000100100110;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1000100100010;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1000100011110;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1000100011001;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1000100010101;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1000100010001;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1000100001100;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1000100001000;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1000100000100;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1000100000000;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1000011111011;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1000011110111;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1000011110011;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1000011101111;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000: n6154 = 13'b1000011101010;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000: n6154 = 13'b1000011100110;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000: n6154 = 13'b1000011100010;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000: n6154 = 13'b1000011011110;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000: n6154 = 13'b1000011011010;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000: n6154 = 13'b1000011010101;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000: n6154 = 13'b1000011010001;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000: n6154 = 13'b1000011001101;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000: n6154 = 13'b1000011001001;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000: n6154 = 13'b1000011000101;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000: n6154 = 13'b1000011000000;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000: n6154 = 13'b1000010111100;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000: n6154 = 13'b1000010111000;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000: n6154 = 13'b1000010110100;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000: n6154 = 13'b1000010110000;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000: n6154 = 13'b1000010101011;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000: n6154 = 13'b1000010100111;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000: n6154 = 13'b1000010100011;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000: n6154 = 13'b1000010011111;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000: n6154 = 13'b1000010011011;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000: n6154 = 13'b1000010010111;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000: n6154 = 13'b1000010010011;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000: n6154 = 13'b1000010001110;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000: n6154 = 13'b1000010001010;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000: n6154 = 13'b1000010000110;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000: n6154 = 13'b1000010000010;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000: n6154 = 13'b1000001111110;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000: n6154 = 13'b1000001111010;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000: n6154 = 13'b1000001110110;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000: n6154 = 13'b1000001110010;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000: n6154 = 13'b1000001101101;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000: n6154 = 13'b1000001101001;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000: n6154 = 13'b1000001100101;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000: n6154 = 13'b1000001100001;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000: n6154 = 13'b1000001011101;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000: n6154 = 13'b1000001011001;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000: n6154 = 13'b1000001010101;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000: n6154 = 13'b1000001010001;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000: n6154 = 13'b1000001001101;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000: n6154 = 13'b1000001001001;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000: n6154 = 13'b1000001000101;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000: n6154 = 13'b1000001000001;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000: n6154 = 13'b1000000111100;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000: n6154 = 13'b1000000111000;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000: n6154 = 13'b1000000110100;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000: n6154 = 13'b1000000110000;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000: n6154 = 13'b1000000101100;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000: n6154 = 13'b1000000101000;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000: n6154 = 13'b1000000100100;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000: n6154 = 13'b1000000100000;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000: n6154 = 13'b1000000011100;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000: n6154 = 13'b1000000011000;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000: n6154 = 13'b1000000010100;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000: n6154 = 13'b1000000010000;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000: n6154 = 13'b1000000001100;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100: n6154 = 13'b1000000001000;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010: n6154 = 13'b1000000000100;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001: n6154 = 13'b1000000000000;
      default: n6154 = 13'bX;
    endcase
endmodule

module intadder_10_freq500_uid102
  (input  clk,
   input  [9:0] x,
   input  [9:0] y,
   input  cin,
   output [9:0] r);
  wire [9:0] rtmp;
  wire [9:0] x_d1;
  wire [9:0] x_d2;
  wire cin_d1;
  wire cin_d2;
  wire cin_d3;
  wire cin_d4;
  wire cin_d5;
  wire cin_d6;
  wire cin_d7;
  wire cin_d8;
  wire cin_d9;
  wire cin_d10;
  wire cin_d11;
  wire cin_d12;
  wire cin_d13;
  wire cin_d14;
  wire cin_d15;
  wire cin_d16;
  wire cin_d17;
  wire [9:0] n3057;
  wire [9:0] n3058;
  wire [9:0] n3059;
  reg [9:0] n3060;
  reg [9:0] n3061;
  reg n3062;
  reg n3063;
  reg n3064;
  reg n3065;
  reg n3066;
  reg n3067;
  reg n3068;
  reg n3069;
  reg n3070;
  reg n3071;
  reg n3072;
  reg n3073;
  reg n3074;
  reg n3075;
  reg n3076;
  reg n3077;
  reg n3078;
  assign r = rtmp; //(module output)
  /* fppowbf16.vhdl:4565:8  */
  assign rtmp = n3059; // (signal)
  /* fppowbf16.vhdl:4567:8  */
  assign x_d1 = n3060; // (signal)
  /* fppowbf16.vhdl:4567:14  */
  assign x_d2 = n3061; // (signal)
  /* fppowbf16.vhdl:4569:8  */
  assign cin_d1 = n3062; // (signal)
  /* fppowbf16.vhdl:4569:16  */
  assign cin_d2 = n3063; // (signal)
  /* fppowbf16.vhdl:4569:24  */
  assign cin_d3 = n3064; // (signal)
  /* fppowbf16.vhdl:4569:32  */
  assign cin_d4 = n3065; // (signal)
  /* fppowbf16.vhdl:4569:40  */
  assign cin_d5 = n3066; // (signal)
  /* fppowbf16.vhdl:4569:48  */
  assign cin_d6 = n3067; // (signal)
  /* fppowbf16.vhdl:4569:56  */
  assign cin_d7 = n3068; // (signal)
  /* fppowbf16.vhdl:4569:64  */
  assign cin_d8 = n3069; // (signal)
  /* fppowbf16.vhdl:4569:72  */
  assign cin_d9 = n3070; // (signal)
  /* fppowbf16.vhdl:4569:80  */
  assign cin_d10 = n3071; // (signal)
  /* fppowbf16.vhdl:4569:89  */
  assign cin_d11 = n3072; // (signal)
  /* fppowbf16.vhdl:4569:98  */
  assign cin_d12 = n3073; // (signal)
  /* fppowbf16.vhdl:4569:107  */
  assign cin_d13 = n3074; // (signal)
  /* fppowbf16.vhdl:4569:116  */
  assign cin_d14 = n3075; // (signal)
  /* fppowbf16.vhdl:4569:125  */
  assign cin_d15 = n3076; // (signal)
  /* fppowbf16.vhdl:4569:134  */
  assign cin_d16 = n3077; // (signal)
  /* fppowbf16.vhdl:4569:143  */
  assign cin_d17 = n3078; // (signal)
  /* fppowbf16.vhdl:4596:17  */
  assign n3057 = x_d2 + y;
  /* fppowbf16.vhdl:4596:21  */
  assign n3058 = {9'b0, cin_d17};  //  uext
  /* fppowbf16.vhdl:4596:21  */
  assign n3059 = n3057 + n3058;
  /* fppowbf16.vhdl:4574:10  */
  always @(posedge clk)
    n3060 <= x;
  /* fppowbf16.vhdl:4574:10  */
  always @(posedge clk)
    n3061 <= x_d1;
  /* fppowbf16.vhdl:4574:10  */
  always @(posedge clk)
    n3062 <= cin;
  /* fppowbf16.vhdl:4574:10  */
  always @(posedge clk)
    n3063 <= cin_d1;
  /* fppowbf16.vhdl:4574:10  */
  always @(posedge clk)
    n3064 <= cin_d2;
  /* fppowbf16.vhdl:4574:10  */
  always @(posedge clk)
    n3065 <= cin_d3;
  /* fppowbf16.vhdl:4574:10  */
  always @(posedge clk)
    n3066 <= cin_d4;
  /* fppowbf16.vhdl:4574:10  */
  always @(posedge clk)
    n3067 <= cin_d5;
  /* fppowbf16.vhdl:4574:10  */
  always @(posedge clk)
    n3068 <= cin_d6;
  /* fppowbf16.vhdl:4574:10  */
  always @(posedge clk)
    n3069 <= cin_d7;
  /* fppowbf16.vhdl:4574:10  */
  always @(posedge clk)
    n3070 <= cin_d8;
  /* fppowbf16.vhdl:4574:10  */
  always @(posedge clk)
    n3071 <= cin_d9;
  /* fppowbf16.vhdl:4574:10  */
  always @(posedge clk)
    n3072 <= cin_d10;
  /* fppowbf16.vhdl:4574:10  */
  always @(posedge clk)
    n3073 <= cin_d11;
  /* fppowbf16.vhdl:4574:10  */
  always @(posedge clk)
    n3074 <= cin_d12;
  /* fppowbf16.vhdl:4574:10  */
  always @(posedge clk)
    n3075 <= cin_d13;
  /* fppowbf16.vhdl:4574:10  */
  always @(posedge clk)
    n3076 <= cin_d14;
  /* fppowbf16.vhdl:4574:10  */
  always @(posedge clk)
    n3077 <= cin_d15;
  /* fppowbf16.vhdl:4574:10  */
  always @(posedge clk)
    n3078 <= cin_d16;
endmodule

module fixrealkcm_freq500_uid89
  (input  clk,
   input  [7:0] x,
   output [17:0] r);
  wire [4:0] fixrealkcm_freq500_uid89_a0;
  wire [17:0] fixrealkcm_freq500_uid89_t0;
  wire [17:0] fixrealkcm_freq500_uid89_t0_copy93;
  wire bh90_w0_0;
  wire bh90_w1_0;
  wire bh90_w2_0;
  wire bh90_w3_0;
  wire bh90_w4_0;
  wire bh90_w5_0;
  wire bh90_w6_0;
  wire bh90_w7_0;
  wire bh90_w8_0;
  wire bh90_w9_0;
  wire bh90_w10_0;
  wire bh90_w11_0;
  wire bh90_w12_0;
  wire bh90_w13_0;
  wire bh90_w14_0;
  wire bh90_w15_0;
  wire bh90_w16_0;
  wire bh90_w17_0;
  wire [2:0] fixrealkcm_freq500_uid89_a1;
  wire [12:0] fixrealkcm_freq500_uid89_t1;
  wire [12:0] fixrealkcm_freq500_uid89_t1_copy96;
  wire bh90_w0_1;
  wire bh90_w1_1;
  wire bh90_w2_1;
  wire bh90_w3_1;
  wire bh90_w4_1;
  wire bh90_w5_1;
  wire bh90_w6_1;
  wire bh90_w7_1;
  wire bh90_w8_1;
  wire bh90_w9_1;
  wire bh90_w10_1;
  wire bh90_w11_1;
  wire bh90_w12_1;
  wire [17:0] bitheapfinaladd_bh90_in0;
  wire [17:0] bitheapfinaladd_bh90_in1;
  wire bitheapfinaladd_bh90_cin;
  wire [17:0] bitheapfinaladd_bh90_out;
  wire [17:0] bitheapresult_bh90;
  wire [17:0] outres;
  wire [4:0] n2958;
  wire [17:0] fixrealkcm_freq500_uid89_table0_n2959;
  wire n2962;
  wire n2963;
  wire n2964;
  wire n2965;
  wire n2966;
  wire n2967;
  wire n2968;
  wire n2969;
  wire n2970;
  wire n2971;
  wire n2972;
  wire n2973;
  wire n2974;
  wire n2975;
  wire n2976;
  wire n2977;
  wire n2978;
  wire n2979;
  wire [2:0] n2980;
  wire [12:0] fixrealkcm_freq500_uid89_table1_n2981;
  wire n2984;
  wire n2985;
  wire n2986;
  wire n2987;
  wire n2988;
  wire n2989;
  wire n2990;
  wire n2991;
  wire n2992;
  wire n2993;
  wire n2994;
  wire n2995;
  wire n2996;
  wire [1:0] n2998;
  wire [2:0] n2999;
  wire [3:0] n3000;
  wire [4:0] n3001;
  wire [5:0] n3002;
  wire [6:0] n3003;
  wire [7:0] n3004;
  wire [8:0] n3005;
  wire [9:0] n3006;
  wire [10:0] n3007;
  wire [11:0] n3008;
  wire [12:0] n3009;
  wire [13:0] n3010;
  wire [14:0] n3011;
  wire [15:0] n3012;
  wire [16:0] n3013;
  wire [17:0] n3014;
  wire [5:0] n3016;
  wire [6:0] n3017;
  wire [7:0] n3018;
  wire [8:0] n3019;
  wire [9:0] n3020;
  wire [10:0] n3021;
  wire [11:0] n3022;
  wire [12:0] n3023;
  wire [13:0] n3024;
  wire [14:0] n3025;
  wire [15:0] n3026;
  wire [16:0] n3027;
  wire [17:0] n3028;
  wire [17:0] bitheapfinaladd_bh90_n3030;
  assign r = outres; //(module output)
  /* fppowbf16.vhdl:4384:8  */
  assign fixrealkcm_freq500_uid89_a0 = n2958; // (signal)
  /* fppowbf16.vhdl:4386:8  */
  assign fixrealkcm_freq500_uid89_t0 = fixrealkcm_freq500_uid89_t0_copy93; // (signal)
  /* fppowbf16.vhdl:4388:8  */
  assign fixrealkcm_freq500_uid89_t0_copy93 = fixrealkcm_freq500_uid89_table0_n2959; // (signal)
  /* fppowbf16.vhdl:4390:8  */
  assign bh90_w0_0 = n2962; // (signal)
  /* fppowbf16.vhdl:4392:8  */
  assign bh90_w1_0 = n2963; // (signal)
  /* fppowbf16.vhdl:4394:8  */
  assign bh90_w2_0 = n2964; // (signal)
  /* fppowbf16.vhdl:4396:8  */
  assign bh90_w3_0 = n2965; // (signal)
  /* fppowbf16.vhdl:4398:8  */
  assign bh90_w4_0 = n2966; // (signal)
  /* fppowbf16.vhdl:4400:8  */
  assign bh90_w5_0 = n2967; // (signal)
  /* fppowbf16.vhdl:4402:8  */
  assign bh90_w6_0 = n2968; // (signal)
  /* fppowbf16.vhdl:4404:8  */
  assign bh90_w7_0 = n2969; // (signal)
  /* fppowbf16.vhdl:4406:8  */
  assign bh90_w8_0 = n2970; // (signal)
  /* fppowbf16.vhdl:4408:8  */
  assign bh90_w9_0 = n2971; // (signal)
  /* fppowbf16.vhdl:4410:8  */
  assign bh90_w10_0 = n2972; // (signal)
  /* fppowbf16.vhdl:4412:8  */
  assign bh90_w11_0 = n2973; // (signal)
  /* fppowbf16.vhdl:4414:8  */
  assign bh90_w12_0 = n2974; // (signal)
  /* fppowbf16.vhdl:4416:8  */
  assign bh90_w13_0 = n2975; // (signal)
  /* fppowbf16.vhdl:4418:8  */
  assign bh90_w14_0 = n2976; // (signal)
  /* fppowbf16.vhdl:4420:8  */
  assign bh90_w15_0 = n2977; // (signal)
  /* fppowbf16.vhdl:4422:8  */
  assign bh90_w16_0 = n2978; // (signal)
  /* fppowbf16.vhdl:4518:35  */
  assign bh90_w17_0 = n2979; // (signal)
  /* fppowbf16.vhdl:4426:8  */
  assign fixrealkcm_freq500_uid89_a1 = n2980; // (signal)
  /* fppowbf16.vhdl:4428:8  */
  assign fixrealkcm_freq500_uid89_t1 = fixrealkcm_freq500_uid89_t1_copy96; // (signal)
  /* fppowbf16.vhdl:4430:8  */
  assign fixrealkcm_freq500_uid89_t1_copy96 = fixrealkcm_freq500_uid89_table1_n2981; // (signal)
  /* fppowbf16.vhdl:4432:8  */
  assign bh90_w0_1 = n2984; // (signal)
  /* fppowbf16.vhdl:4434:8  */
  assign bh90_w1_1 = n2985; // (signal)
  /* fppowbf16.vhdl:4436:8  */
  assign bh90_w2_1 = n2986; // (signal)
  /* fppowbf16.vhdl:4438:8  */
  assign bh90_w3_1 = n2987; // (signal)
  /* fppowbf16.vhdl:4440:8  */
  assign bh90_w4_1 = n2988; // (signal)
  /* fppowbf16.vhdl:4442:8  */
  assign bh90_w5_1 = n2989; // (signal)
  /* fppowbf16.vhdl:4444:8  */
  assign bh90_w6_1 = n2990; // (signal)
  /* fppowbf16.vhdl:4446:8  */
  assign bh90_w7_1 = n2991; // (signal)
  /* fppowbf16.vhdl:4448:8  */
  assign bh90_w8_1 = n2992; // (signal)
  /* fppowbf16.vhdl:4450:8  */
  assign bh90_w9_1 = n2993; // (signal)
  /* fppowbf16.vhdl:4452:8  */
  assign bh90_w10_1 = n2994; // (signal)
  /* fppowbf16.vhdl:4454:8  */
  assign bh90_w11_1 = n2995; // (signal)
  /* fppowbf16.vhdl:4456:8  */
  assign bh90_w12_1 = n2996; // (signal)
  /* fppowbf16.vhdl:4458:8  */
  assign bitheapfinaladd_bh90_in0 = n3014; // (signal)
  /* fppowbf16.vhdl:4460:8  */
  assign bitheapfinaladd_bh90_in1 = n3028; // (signal)
  /* fppowbf16.vhdl:4462:8  */
  assign bitheapfinaladd_bh90_cin = 1'b0; // (signal)
  /* fppowbf16.vhdl:4464:8  */
  assign bitheapfinaladd_bh90_out = bitheapfinaladd_bh90_n3030; // (signal)
  /* fppowbf16.vhdl:4466:8  */
  assign bitheapresult_bh90 = bitheapfinaladd_bh90_out; // (signal)
  /* fppowbf16.vhdl:4468:8  */
  assign outres = bitheapresult_bh90; // (signal)
  /* fppowbf16.vhdl:4472:36  */
  assign n2958 = x[7:3]; // extract
  /* fppowbf16.vhdl:4473:4  */
  fixrealkcm_freq500_uid89_t0_freq500_uid92 fixrealkcm_freq500_uid89_table0 (
    .x(fixrealkcm_freq500_uid89_a0),
    .y(fixrealkcm_freq500_uid89_table0_n2959));
  /* fppowbf16.vhdl:4477:44  */
  assign n2962 = fixrealkcm_freq500_uid89_t0[0]; // extract
  /* fppowbf16.vhdl:4478:44  */
  assign n2963 = fixrealkcm_freq500_uid89_t0[1]; // extract
  /* fppowbf16.vhdl:4479:44  */
  assign n2964 = fixrealkcm_freq500_uid89_t0[2]; // extract
  /* fppowbf16.vhdl:4480:44  */
  assign n2965 = fixrealkcm_freq500_uid89_t0[3]; // extract
  /* fppowbf16.vhdl:4481:44  */
  assign n2966 = fixrealkcm_freq500_uid89_t0[4]; // extract
  /* fppowbf16.vhdl:4482:44  */
  assign n2967 = fixrealkcm_freq500_uid89_t0[5]; // extract
  /* fppowbf16.vhdl:4483:44  */
  assign n2968 = fixrealkcm_freq500_uid89_t0[6]; // extract
  /* fppowbf16.vhdl:4484:44  */
  assign n2969 = fixrealkcm_freq500_uid89_t0[7]; // extract
  /* fppowbf16.vhdl:4485:44  */
  assign n2970 = fixrealkcm_freq500_uid89_t0[8]; // extract
  /* fppowbf16.vhdl:4486:44  */
  assign n2971 = fixrealkcm_freq500_uid89_t0[9]; // extract
  /* fppowbf16.vhdl:4487:45  */
  assign n2972 = fixrealkcm_freq500_uid89_t0[10]; // extract
  /* fppowbf16.vhdl:4488:45  */
  assign n2973 = fixrealkcm_freq500_uid89_t0[11]; // extract
  /* fppowbf16.vhdl:4489:45  */
  assign n2974 = fixrealkcm_freq500_uid89_t0[12]; // extract
  /* fppowbf16.vhdl:4490:45  */
  assign n2975 = fixrealkcm_freq500_uid89_t0[13]; // extract
  /* fppowbf16.vhdl:4491:45  */
  assign n2976 = fixrealkcm_freq500_uid89_t0[14]; // extract
  /* fppowbf16.vhdl:4492:45  */
  assign n2977 = fixrealkcm_freq500_uid89_t0[15]; // extract
  /* fppowbf16.vhdl:4493:45  */
  assign n2978 = fixrealkcm_freq500_uid89_t0[16]; // extract
  /* fppowbf16.vhdl:4494:45  */
  assign n2979 = fixrealkcm_freq500_uid89_t0[17]; // extract
  /* fppowbf16.vhdl:4495:36  */
  assign n2980 = x[2:0]; // extract
  /* fppowbf16.vhdl:4496:4  */
  fixrealkcm_freq500_uid89_t1_freq500_uid95 fixrealkcm_freq500_uid89_table1 (
    .x(fixrealkcm_freq500_uid89_a1),
    .y(fixrealkcm_freq500_uid89_table1_n2981));
  /* fppowbf16.vhdl:4500:44  */
  assign n2984 = fixrealkcm_freq500_uid89_t1[0]; // extract
  /* fppowbf16.vhdl:4501:44  */
  assign n2985 = fixrealkcm_freq500_uid89_t1[1]; // extract
  /* fppowbf16.vhdl:4502:44  */
  assign n2986 = fixrealkcm_freq500_uid89_t1[2]; // extract
  /* fppowbf16.vhdl:4503:44  */
  assign n2987 = fixrealkcm_freq500_uid89_t1[3]; // extract
  /* fppowbf16.vhdl:4504:44  */
  assign n2988 = fixrealkcm_freq500_uid89_t1[4]; // extract
  /* fppowbf16.vhdl:4505:44  */
  assign n2989 = fixrealkcm_freq500_uid89_t1[5]; // extract
  /* fppowbf16.vhdl:4506:44  */
  assign n2990 = fixrealkcm_freq500_uid89_t1[6]; // extract
  /* fppowbf16.vhdl:4507:44  */
  assign n2991 = fixrealkcm_freq500_uid89_t1[7]; // extract
  /* fppowbf16.vhdl:4508:44  */
  assign n2992 = fixrealkcm_freq500_uid89_t1[8]; // extract
  /* fppowbf16.vhdl:4509:44  */
  assign n2993 = fixrealkcm_freq500_uid89_t1[9]; // extract
  /* fppowbf16.vhdl:4510:45  */
  assign n2994 = fixrealkcm_freq500_uid89_t1[10]; // extract
  /* fppowbf16.vhdl:4511:45  */
  assign n2995 = fixrealkcm_freq500_uid89_t1[11]; // extract
  /* fppowbf16.vhdl:4512:45  */
  assign n2996 = fixrealkcm_freq500_uid89_t1[12]; // extract
  /* fppowbf16.vhdl:4518:48  */
  assign n2998 = {bh90_w17_0, bh90_w16_0};
  /* fppowbf16.vhdl:4518:61  */
  assign n2999 = {n2998, bh90_w15_0};
  /* fppowbf16.vhdl:4518:74  */
  assign n3000 = {n2999, bh90_w14_0};
  /* fppowbf16.vhdl:4518:87  */
  assign n3001 = {n3000, bh90_w13_0};
  /* fppowbf16.vhdl:4518:100  */
  assign n3002 = {n3001, bh90_w12_0};
  /* fppowbf16.vhdl:4518:113  */
  assign n3003 = {n3002, bh90_w11_0};
  /* fppowbf16.vhdl:4518:126  */
  assign n3004 = {n3003, bh90_w10_0};
  /* fppowbf16.vhdl:4518:139  */
  assign n3005 = {n3004, bh90_w9_0};
  /* fppowbf16.vhdl:4518:151  */
  assign n3006 = {n3005, bh90_w8_0};
  /* fppowbf16.vhdl:4518:163  */
  assign n3007 = {n3006, bh90_w7_0};
  /* fppowbf16.vhdl:4518:175  */
  assign n3008 = {n3007, bh90_w6_0};
  /* fppowbf16.vhdl:4518:187  */
  assign n3009 = {n3008, bh90_w5_0};
  /* fppowbf16.vhdl:4518:199  */
  assign n3010 = {n3009, bh90_w4_0};
  /* fppowbf16.vhdl:4518:211  */
  assign n3011 = {n3010, bh90_w3_0};
  /* fppowbf16.vhdl:4518:223  */
  assign n3012 = {n3011, bh90_w2_0};
  /* fppowbf16.vhdl:4518:235  */
  assign n3013 = {n3012, bh90_w1_0};
  /* fppowbf16.vhdl:4518:247  */
  assign n3014 = {n3013, bh90_w0_0};
  /* fppowbf16.vhdl:4519:60  */
  assign n3016 = {5'b00000, bh90_w12_1};
  /* fppowbf16.vhdl:4519:73  */
  assign n3017 = {n3016, bh90_w11_1};
  /* fppowbf16.vhdl:4519:86  */
  assign n3018 = {n3017, bh90_w10_1};
  /* fppowbf16.vhdl:4519:99  */
  assign n3019 = {n3018, bh90_w9_1};
  /* fppowbf16.vhdl:4519:111  */
  assign n3020 = {n3019, bh90_w8_1};
  /* fppowbf16.vhdl:4519:123  */
  assign n3021 = {n3020, bh90_w7_1};
  /* fppowbf16.vhdl:4519:135  */
  assign n3022 = {n3021, bh90_w6_1};
  /* fppowbf16.vhdl:4519:147  */
  assign n3023 = {n3022, bh90_w5_1};
  /* fppowbf16.vhdl:4519:159  */
  assign n3024 = {n3023, bh90_w4_1};
  /* fppowbf16.vhdl:4519:171  */
  assign n3025 = {n3024, bh90_w3_1};
  /* fppowbf16.vhdl:4519:183  */
  assign n3026 = {n3025, bh90_w2_1};
  /* fppowbf16.vhdl:4519:195  */
  assign n3027 = {n3026, bh90_w1_1};
  /* fppowbf16.vhdl:4519:207  */
  assign n3028 = {n3027, bh90_w0_1};
  /* fppowbf16.vhdl:4522:4  */
  intadder_18_freq500_uid99 bitheapfinaladd_bh90 (
    .clk(clk),
    .x(bitheapfinaladd_bh90_in0),
    .y(bitheapfinaladd_bh90_in1),
    .cin(bitheapfinaladd_bh90_cin),
    .r(bitheapfinaladd_bh90_n3030));
endmodule

module fixrealkcm_freq500_uid77
  (input  clk,
   input  [9:0] x,
   output [7:0] r);
  wire [4:0] fixrealkcm_freq500_uid77_a0;
  wire [11:0] fixrealkcm_freq500_uid77_t0;
  wire [11:0] fixrealkcm_freq500_uid77_t0_copy81;
  wire bh78_w0_0;
  wire bh78_w1_0;
  wire bh78_w2_0;
  wire bh78_w3_0;
  wire bh78_w4_0;
  wire bh78_w5_0;
  wire bh78_w6_0;
  wire bh78_w7_0;
  wire bh78_w8_0;
  wire bh78_w9_0;
  wire bh78_w10_0;
  wire bh78_w11_0;
  wire [4:0] fixrealkcm_freq500_uid77_a1;
  wire [6:0] fixrealkcm_freq500_uid77_t1;
  wire [6:0] fixrealkcm_freq500_uid77_t1_copy84;
  wire bh78_w0_1;
  wire bh78_w1_1;
  wire bh78_w2_1;
  wire bh78_w3_1;
  wire bh78_w4_1;
  wire bh78_w5_1;
  wire bh78_w6_1;
  wire [11:0] bitheapfinaladd_bh78_in0;
  wire [11:0] bitheapfinaladd_bh78_in1;
  wire bitheapfinaladd_bh78_cin;
  wire [11:0] bitheapfinaladd_bh78_out;
  wire [11:0] bitheapresult_bh78;
  wire [11:0] outres;
  wire [4:0] n2905;
  wire [11:0] fixrealkcm_freq500_uid77_table0_n2906;
  wire n2909;
  wire n2910;
  wire n2911;
  wire n2912;
  wire n2913;
  wire n2914;
  wire n2915;
  wire n2916;
  wire n2917;
  wire n2918;
  wire n2919;
  wire n2920;
  wire [4:0] n2921;
  wire [6:0] fixrealkcm_freq500_uid77_table1_n2922;
  wire n2925;
  wire n2926;
  wire n2927;
  wire n2928;
  wire n2929;
  wire n2930;
  wire n2931;
  wire [1:0] n2933;
  wire [2:0] n2934;
  wire [3:0] n2935;
  wire [4:0] n2936;
  wire [5:0] n2937;
  wire [6:0] n2938;
  wire [7:0] n2939;
  wire [8:0] n2940;
  wire [9:0] n2941;
  wire [10:0] n2942;
  wire [11:0] n2943;
  wire [5:0] n2945;
  wire [6:0] n2946;
  wire [7:0] n2947;
  wire [8:0] n2948;
  wire [9:0] n2949;
  wire [10:0] n2950;
  wire [11:0] n2951;
  wire [11:0] bitheapfinaladd_bh78_n2953;
  wire [7:0] n2956;
  assign r = n2956; //(module output)
  /* fppowbf16.vhdl:4154:8  */
  assign fixrealkcm_freq500_uid77_a0 = n2905; // (signal)
  /* fppowbf16.vhdl:4156:8  */
  assign fixrealkcm_freq500_uid77_t0 = fixrealkcm_freq500_uid77_t0_copy81; // (signal)
  /* fppowbf16.vhdl:4158:8  */
  assign fixrealkcm_freq500_uid77_t0_copy81 = fixrealkcm_freq500_uid77_table0_n2906; // (signal)
  /* fppowbf16.vhdl:4160:8  */
  assign bh78_w0_0 = n2909; // (signal)
  /* fppowbf16.vhdl:4162:8  */
  assign bh78_w1_0 = n2910; // (signal)
  /* fppowbf16.vhdl:4164:8  */
  assign bh78_w2_0 = n2911; // (signal)
  /* fppowbf16.vhdl:4166:8  */
  assign bh78_w3_0 = n2912; // (signal)
  /* fppowbf16.vhdl:4168:8  */
  assign bh78_w4_0 = n2913; // (signal)
  /* fppowbf16.vhdl:4170:8  */
  assign bh78_w5_0 = n2914; // (signal)
  /* fppowbf16.vhdl:4172:8  */
  assign bh78_w6_0 = n2915; // (signal)
  /* fppowbf16.vhdl:4174:8  */
  assign bh78_w7_0 = n2916; // (signal)
  /* fppowbf16.vhdl:4176:8  */
  assign bh78_w8_0 = n2917; // (signal)
  /* fppowbf16.vhdl:4178:8  */
  assign bh78_w9_0 = n2918; // (signal)
  /* fppowbf16.vhdl:4180:8  */
  assign bh78_w10_0 = n2919; // (signal)
  /* fppowbf16.vhdl:4252:35  */
  assign bh78_w11_0 = n2920; // (signal)
  /* fppowbf16.vhdl:4184:8  */
  assign fixrealkcm_freq500_uid77_a1 = n2921; // (signal)
  /* fppowbf16.vhdl:4186:8  */
  assign fixrealkcm_freq500_uid77_t1 = fixrealkcm_freq500_uid77_t1_copy84; // (signal)
  /* fppowbf16.vhdl:4188:8  */
  assign fixrealkcm_freq500_uid77_t1_copy84 = fixrealkcm_freq500_uid77_table1_n2922; // (signal)
  /* fppowbf16.vhdl:4190:8  */
  assign bh78_w0_1 = n2925; // (signal)
  /* fppowbf16.vhdl:4192:8  */
  assign bh78_w1_1 = n2926; // (signal)
  /* fppowbf16.vhdl:4194:8  */
  assign bh78_w2_1 = n2927; // (signal)
  /* fppowbf16.vhdl:4196:8  */
  assign bh78_w3_1 = n2928; // (signal)
  /* fppowbf16.vhdl:4198:8  */
  assign bh78_w4_1 = n2929; // (signal)
  /* fppowbf16.vhdl:4200:8  */
  assign bh78_w5_1 = n2930; // (signal)
  /* fppowbf16.vhdl:4202:8  */
  assign bh78_w6_1 = n2931; // (signal)
  /* fppowbf16.vhdl:4204:8  */
  assign bitheapfinaladd_bh78_in0 = n2943; // (signal)
  /* fppowbf16.vhdl:4206:8  */
  assign bitheapfinaladd_bh78_in1 = n2951; // (signal)
  /* fppowbf16.vhdl:4208:8  */
  assign bitheapfinaladd_bh78_cin = 1'b0; // (signal)
  /* fppowbf16.vhdl:4210:8  */
  assign bitheapfinaladd_bh78_out = bitheapfinaladd_bh78_n2953; // (signal)
  /* fppowbf16.vhdl:4212:8  */
  assign bitheapresult_bh78 = bitheapfinaladd_bh78_out; // (signal)
  /* fppowbf16.vhdl:4214:8  */
  assign outres = bitheapresult_bh78; // (signal)
  /* fppowbf16.vhdl:4218:36  */
  assign n2905 = x[9:5]; // extract
  /* fppowbf16.vhdl:4219:4  */
  fixrealkcm_freq500_uid77_t0_freq500_uid80 fixrealkcm_freq500_uid77_table0 (
    .x(fixrealkcm_freq500_uid77_a0),
    .y(fixrealkcm_freq500_uid77_table0_n2906));
  /* fppowbf16.vhdl:4223:44  */
  assign n2909 = fixrealkcm_freq500_uid77_t0[0]; // extract
  /* fppowbf16.vhdl:4224:44  */
  assign n2910 = fixrealkcm_freq500_uid77_t0[1]; // extract
  /* fppowbf16.vhdl:4225:44  */
  assign n2911 = fixrealkcm_freq500_uid77_t0[2]; // extract
  /* fppowbf16.vhdl:4226:44  */
  assign n2912 = fixrealkcm_freq500_uid77_t0[3]; // extract
  /* fppowbf16.vhdl:4227:44  */
  assign n2913 = fixrealkcm_freq500_uid77_t0[4]; // extract
  /* fppowbf16.vhdl:4228:44  */
  assign n2914 = fixrealkcm_freq500_uid77_t0[5]; // extract
  /* fppowbf16.vhdl:4229:44  */
  assign n2915 = fixrealkcm_freq500_uid77_t0[6]; // extract
  /* fppowbf16.vhdl:4230:44  */
  assign n2916 = fixrealkcm_freq500_uid77_t0[7]; // extract
  /* fppowbf16.vhdl:4231:44  */
  assign n2917 = fixrealkcm_freq500_uid77_t0[8]; // extract
  /* fppowbf16.vhdl:4232:44  */
  assign n2918 = fixrealkcm_freq500_uid77_t0[9]; // extract
  /* fppowbf16.vhdl:4233:45  */
  assign n2919 = fixrealkcm_freq500_uid77_t0[10]; // extract
  /* fppowbf16.vhdl:4234:45  */
  assign n2920 = fixrealkcm_freq500_uid77_t0[11]; // extract
  /* fppowbf16.vhdl:4235:36  */
  assign n2921 = x[4:0]; // extract
  /* fppowbf16.vhdl:4236:4  */
  fixrealkcm_freq500_uid77_t1_freq500_uid83 fixrealkcm_freq500_uid77_table1 (
    .x(fixrealkcm_freq500_uid77_a1),
    .y(fixrealkcm_freq500_uid77_table1_n2922));
  /* fppowbf16.vhdl:4240:44  */
  assign n2925 = fixrealkcm_freq500_uid77_t1[0]; // extract
  /* fppowbf16.vhdl:4241:44  */
  assign n2926 = fixrealkcm_freq500_uid77_t1[1]; // extract
  /* fppowbf16.vhdl:4242:44  */
  assign n2927 = fixrealkcm_freq500_uid77_t1[2]; // extract
  /* fppowbf16.vhdl:4243:44  */
  assign n2928 = fixrealkcm_freq500_uid77_t1[3]; // extract
  /* fppowbf16.vhdl:4244:44  */
  assign n2929 = fixrealkcm_freq500_uid77_t1[4]; // extract
  /* fppowbf16.vhdl:4245:44  */
  assign n2930 = fixrealkcm_freq500_uid77_t1[5]; // extract
  /* fppowbf16.vhdl:4246:44  */
  assign n2931 = fixrealkcm_freq500_uid77_t1[6]; // extract
  /* fppowbf16.vhdl:4252:48  */
  assign n2933 = {bh78_w11_0, bh78_w10_0};
  /* fppowbf16.vhdl:4252:61  */
  assign n2934 = {n2933, bh78_w9_0};
  /* fppowbf16.vhdl:4252:73  */
  assign n2935 = {n2934, bh78_w8_0};
  /* fppowbf16.vhdl:4252:85  */
  assign n2936 = {n2935, bh78_w7_0};
  /* fppowbf16.vhdl:4252:97  */
  assign n2937 = {n2936, bh78_w6_0};
  /* fppowbf16.vhdl:4252:109  */
  assign n2938 = {n2937, bh78_w5_0};
  /* fppowbf16.vhdl:4252:121  */
  assign n2939 = {n2938, bh78_w4_0};
  /* fppowbf16.vhdl:4252:133  */
  assign n2940 = {n2939, bh78_w3_0};
  /* fppowbf16.vhdl:4252:145  */
  assign n2941 = {n2940, bh78_w2_0};
  /* fppowbf16.vhdl:4252:157  */
  assign n2942 = {n2941, bh78_w1_0};
  /* fppowbf16.vhdl:4252:169  */
  assign n2943 = {n2942, bh78_w0_0};
  /* fppowbf16.vhdl:4253:60  */
  assign n2945 = {5'b00000, bh78_w6_1};
  /* fppowbf16.vhdl:4253:72  */
  assign n2946 = {n2945, bh78_w5_1};
  /* fppowbf16.vhdl:4253:84  */
  assign n2947 = {n2946, bh78_w4_1};
  /* fppowbf16.vhdl:4253:96  */
  assign n2948 = {n2947, bh78_w3_1};
  /* fppowbf16.vhdl:4253:108  */
  assign n2949 = {n2948, bh78_w2_1};
  /* fppowbf16.vhdl:4253:120  */
  assign n2950 = {n2949, bh78_w1_1};
  /* fppowbf16.vhdl:4253:132  */
  assign n2951 = {n2950, bh78_w0_1};
  /* fppowbf16.vhdl:4256:4  */
  intadder_12_freq500_uid87 bitheapfinaladd_bh78 (
    .clk(clk),
    .x(bitheapfinaladd_bh78_in0),
    .y(bitheapfinaladd_bh78_in1),
    .cin(bitheapfinaladd_bh78_cin),
    .r(bitheapfinaladd_bh78_n2953));
  /* fppowbf16.vhdl:4264:15  */
  assign n2956 = outres[11:4]; // extract
endmodule

module intadder_29_freq500_uid49
  (input  clk,
   input  [28:0] x,
   input  [28:0] y,
   input  cin,
   output [28:0] r);
  wire [28:0] rtmp;
  wire cin_d1;
  wire [28:0] n2900;
  wire [28:0] n2901;
  wire [28:0] n2902;
  reg n2903;
  assign r = rtmp; //(module output)
  /* fppowbf16.vhdl:2445:8  */
  assign rtmp = n2902; // (signal)
  /* fppowbf16.vhdl:2447:8  */
  assign cin_d1 = n2903; // (signal)
  /* fppowbf16.vhdl:2456:14  */
  assign n2900 = x + y;
  /* fppowbf16.vhdl:2456:18  */
  assign n2901 = {28'b0, cin_d1};  //  uext
  /* fppowbf16.vhdl:2456:18  */
  assign n2902 = n2900 + n2901;
  /* fppowbf16.vhdl:2452:10  */
  always @(posedge clk)
    n2903 <= cin;
endmodule

module fixrealkcm_freq500_uid39_t1_freq500_uid45
  (input  [2:0] x,
   output [23:0] y);
  wire [23:0] y0;
  wire [23:0] y1;
  wire n2869;
  wire n2872;
  wire n2875;
  wire n2878;
  wire n2881;
  wire n2884;
  wire n2887;
  wire n2890;
  wire [7:0] n2892;
  reg [23:0] n2893;
  assign y = y1; //(module output)
  /* fppowbf16.vhdl:510:8  */
  assign y0 = n2893; // (signal)
  /* fppowbf16.vhdl:512:8  */
  assign y1 = y0; // (signal)
  /* fppowbf16.vhdl:516:34  */
  assign n2869 = x == 3'b000;
  /* fppowbf16.vhdl:517:34  */
  assign n2872 = x == 3'b001;
  /* fppowbf16.vhdl:518:34  */
  assign n2875 = x == 3'b010;
  /* fppowbf16.vhdl:519:34  */
  assign n2878 = x == 3'b011;
  /* fppowbf16.vhdl:520:34  */
  assign n2881 = x == 3'b100;
  /* fppowbf16.vhdl:521:34  */
  assign n2884 = x == 3'b101;
  /* fppowbf16.vhdl:522:34  */
  assign n2887 = x == 3'b110;
  /* fppowbf16.vhdl:523:34  */
  assign n2890 = x == 3'b111;
  assign n2892 = {n2890, n2887, n2884, n2881, n2878, n2875, n2872, n2869};
  /* fppowbf16.vhdl:515:4  */
  always @*
    case (n2892)
      8'b10000000: n2893 = 24'b100110110100001111010101;
      8'b01000000: n2893 = 24'b100001010001010110010010;
      8'b00100000: n2893 = 24'b011011101110011101001111;
      8'b00010000: n2893 = 24'b010110001011100100001100;
      8'b00001000: n2893 = 24'b010000101000101011001001;
      8'b00000100: n2893 = 24'b001011000101110010000110;
      8'b00000010: n2893 = 24'b000101100010111001000011;
      8'b00000001: n2893 = 24'b000000000000000000000000;
      default: n2893 = 24'bX;
    endcase
endmodule

module fixrealkcm_freq500_uid39_t0_freq500_uid42
  (input  [4:0] x,
   output [28:0] y);
  wire [28:0] y0;
  wire [28:0] y1;
  wire n2769;
  wire n2772;
  wire n2775;
  wire n2778;
  wire n2781;
  wire n2784;
  wire n2787;
  wire n2790;
  wire n2793;
  wire n2796;
  wire n2799;
  wire n2802;
  wire n2805;
  wire n2808;
  wire n2811;
  wire n2814;
  wire n2817;
  wire n2820;
  wire n2823;
  wire n2826;
  wire n2829;
  wire n2832;
  wire n2835;
  wire n2838;
  wire n2841;
  wire n2844;
  wire n2847;
  wire n2850;
  wire n2853;
  wire n2856;
  wire n2859;
  wire n2862;
  wire [31:0] n2864;
  reg [28:0] n2865;
  assign y = y1; //(module output)
  /* fppowbf16.vhdl:438:8  */
  assign y0 = n2865; // (signal)
  /* fppowbf16.vhdl:440:8  */
  assign y1 = y0; // (signal)
  /* fppowbf16.vhdl:444:39  */
  assign n2769 = x == 5'b00000;
  /* fppowbf16.vhdl:445:39  */
  assign n2772 = x == 5'b00001;
  /* fppowbf16.vhdl:446:39  */
  assign n2775 = x == 5'b00010;
  /* fppowbf16.vhdl:447:39  */
  assign n2778 = x == 5'b00011;
  /* fppowbf16.vhdl:448:39  */
  assign n2781 = x == 5'b00100;
  /* fppowbf16.vhdl:449:39  */
  assign n2784 = x == 5'b00101;
  /* fppowbf16.vhdl:450:39  */
  assign n2787 = x == 5'b00110;
  /* fppowbf16.vhdl:451:39  */
  assign n2790 = x == 5'b00111;
  /* fppowbf16.vhdl:452:39  */
  assign n2793 = x == 5'b01000;
  /* fppowbf16.vhdl:453:39  */
  assign n2796 = x == 5'b01001;
  /* fppowbf16.vhdl:454:39  */
  assign n2799 = x == 5'b01010;
  /* fppowbf16.vhdl:455:39  */
  assign n2802 = x == 5'b01011;
  /* fppowbf16.vhdl:456:39  */
  assign n2805 = x == 5'b01100;
  /* fppowbf16.vhdl:457:39  */
  assign n2808 = x == 5'b01101;
  /* fppowbf16.vhdl:458:39  */
  assign n2811 = x == 5'b01110;
  /* fppowbf16.vhdl:459:39  */
  assign n2814 = x == 5'b01111;
  /* fppowbf16.vhdl:460:39  */
  assign n2817 = x == 5'b10000;
  /* fppowbf16.vhdl:461:39  */
  assign n2820 = x == 5'b10001;
  /* fppowbf16.vhdl:462:39  */
  assign n2823 = x == 5'b10010;
  /* fppowbf16.vhdl:463:39  */
  assign n2826 = x == 5'b10011;
  /* fppowbf16.vhdl:464:39  */
  assign n2829 = x == 5'b10100;
  /* fppowbf16.vhdl:465:39  */
  assign n2832 = x == 5'b10101;
  /* fppowbf16.vhdl:466:39  */
  assign n2835 = x == 5'b10110;
  /* fppowbf16.vhdl:467:39  */
  assign n2838 = x == 5'b10111;
  /* fppowbf16.vhdl:468:39  */
  assign n2841 = x == 5'b11000;
  /* fppowbf16.vhdl:469:39  */
  assign n2844 = x == 5'b11001;
  /* fppowbf16.vhdl:470:39  */
  assign n2847 = x == 5'b11010;
  /* fppowbf16.vhdl:471:39  */
  assign n2850 = x == 5'b11011;
  /* fppowbf16.vhdl:472:39  */
  assign n2853 = x == 5'b11100;
  /* fppowbf16.vhdl:473:39  */
  assign n2856 = x == 5'b11101;
  /* fppowbf16.vhdl:474:39  */
  assign n2859 = x == 5'b11110;
  /* fppowbf16.vhdl:475:39  */
  assign n2862 = x == 5'b11111;
  assign n2864 = {n2862, n2859, n2856, n2853, n2850, n2847, n2844, n2841, n2838, n2835, n2832, n2829, n2826, n2823, n2820, n2817, n2814, n2811, n2808, n2805, n2802, n2799, n2796, n2793, n2790, n2787, n2784, n2781, n2778, n2775, n2772, n2769};
  /* fppowbf16.vhdl:443:4  */
  always @*
    case (n2864)
      32'b10000000000000000000000000000000: n2865 = 29'b10101011111001101000011100111;
      32'b01000000000000000000000000000000: n2865 = 29'b10100110010110101111011001111;
      32'b00100000000000000000000000000000: n2865 = 29'b10100000110011110110010110111;
      32'b00010000000000000000000000000000: n2865 = 29'b10011011010000111101010011111;
      32'b00001000000000000000000000000000: n2865 = 29'b10010101101110000100010000111;
      32'b00000100000000000000000000000000: n2865 = 29'b10010000001011001011001101111;
      32'b00000010000000000000000000000000: n2865 = 29'b10001010101000010010001010111;
      32'b00000001000000000000000000000000: n2865 = 29'b10000101000101011001000111111;
      32'b00000000100000000000000000000000: n2865 = 29'b01111111100010100000000100111;
      32'b00000000010000000000000000000000: n2865 = 29'b01111001111111100111000001111;
      32'b00000000001000000000000000000000: n2865 = 29'b01110100011100101101111110111;
      32'b00000000000100000000000000000000: n2865 = 29'b01101110111001110100111011111;
      32'b00000000000010000000000000000000: n2865 = 29'b01101001010110111011111000111;
      32'b00000000000001000000000000000000: n2865 = 29'b01100011110100000010110101111;
      32'b00000000000000100000000000000000: n2865 = 29'b01011110010001001001110010111;
      32'b00000000000000010000000000000000: n2865 = 29'b01011000101110010000101111111;
      32'b00000000000000001000000000000000: n2865 = 29'b01010011001011010111101101000;
      32'b00000000000000000100000000000000: n2865 = 29'b01001101101000011110101010000;
      32'b00000000000000000010000000000000: n2865 = 29'b01001000000101100101100111000;
      32'b00000000000000000001000000000000: n2865 = 29'b01000010100010101100100100000;
      32'b00000000000000000000100000000000: n2865 = 29'b00111100111111110011100001000;
      32'b00000000000000000000010000000000: n2865 = 29'b00110111011100111010011110000;
      32'b00000000000000000000001000000000: n2865 = 29'b00110001111010000001011011000;
      32'b00000000000000000000000100000000: n2865 = 29'b00101100010111001000011000000;
      32'b00000000000000000000000010000000: n2865 = 29'b00100110110100001111010101000;
      32'b00000000000000000000000001000000: n2865 = 29'b00100001010001010110010010000;
      32'b00000000000000000000000000100000: n2865 = 29'b00011011101110011101001111000;
      32'b00000000000000000000000000010000: n2865 = 29'b00010110001011100100001100000;
      32'b00000000000000000000000000001000: n2865 = 29'b00010000101000101011001001000;
      32'b00000000000000000000000000000100: n2865 = 29'b00001011000101110010000110000;
      32'b00000000000000000000000000000010: n2865 = 29'b00000101100010111001000011000;
      32'b00000000000000000000000000000001: n2865 = 29'b00000000000000000000000000000;
      default: n2865 = 29'bX;
    endcase
endmodule

module intadder_17_freq500_uid107
  (input  clk,
   input  [16:0] x,
   input  [16:0] y,
   input  cin,
   output [16:0] r);
  wire [16:0] rtmp;
  wire [16:0] n2763;
  wire [16:0] n2764;
  wire [16:0] n2765;
  assign r = rtmp; //(module output)
  /* fppowbf16.vhdl:4747:8  */
  assign rtmp = n2765; // (signal)
  /* fppowbf16.vhdl:4750:14  */
  assign n2763 = x + y;
  /* fppowbf16.vhdl:4750:18  */
  assign n2764 = {16'b0, cin};  //  uext
  /* fppowbf16.vhdl:4750:18  */
  assign n2765 = n2763 + n2764;
endmodule

module exp_8_7_freq500_uid75
  (input  clk,
   input  [16:0] ufixx_i,
   input  xsign,
   output [12:0] expy,
   output [8:0] k);
  wire [16:0] ufixx;
  wire [9:0] xmulin;
  wire [7:0] absk;
  wire [8:0] minusabsk;
  wire [17:0] absklog2;
  wire [9:0] subop1;
  wire [9:0] subop2;
  wire [9:0] y;
  wire xsign_d1;
  wire xsign_d2;
  wire xsign_d3;
  wire xsign_d4;
  wire [9:0] n2728;
  wire [7:0] mulinvlog2_n2729;
  wire [8:0] n2733;
  wire [8:0] n2735;
  wire [8:0] n2736;
  wire [8:0] n2738;
  wire [17:0] mullog2_n2739;
  wire [9:0] n2742;
  wire n2743;
  wire [9:0] n2744;
  wire [9:0] n2745;
  wire [9:0] n2746;
  wire [9:0] n2747;
  wire [9:0] n2748;
  wire [9:0] n2749;
  wire [9:0] n2750;
  localparam n2751 = 1'b1;
  wire [9:0] theyadder_n2752;
  wire [12:0] expytable_n2755;
  reg n2758;
  reg n2759;
  reg n2760;
  reg n2761;
  assign expy = expytable_n2755; //(module output)
  assign k = n2736; //(module output)
  /* fppowbf16.vhdl:4659:8  */
  assign xmulin = n2728; // (signal)
  /* fppowbf16.vhdl:4661:8  */
  assign absk = mulinvlog2_n2729; // (signal)
  /* fppowbf16.vhdl:4663:8  */
  assign minusabsk = n2735; // (signal)
  /* fppowbf16.vhdl:4665:8  */
  assign absklog2 = mullog2_n2739; // (signal)
  /* fppowbf16.vhdl:4667:8  */
  assign subop1 = n2744; // (signal)
  /* fppowbf16.vhdl:4669:8  */
  assign subop2 = n2748; // (signal)
  /* fppowbf16.vhdl:4671:8  */
  assign y = theyadder_n2752; // (signal)
  /* fppowbf16.vhdl:4673:8  */
  assign xsign_d1 = n2758; // (signal)
  /* fppowbf16.vhdl:4673:18  */
  assign xsign_d2 = n2759; // (signal)
  /* fppowbf16.vhdl:4673:28  */
  assign xsign_d3 = n2760; // (signal)
  /* fppowbf16.vhdl:4673:38  */
  assign xsign_d4 = n2761; // (signal)
  /* fppowbf16.vhdl:4690:19  */
  assign n2728 = ufixx[16:7]; // extract
  /* fppowbf16.vhdl:4691:4  */
  fixrealkcm_freq500_uid77 mulinvlog2 (
    .clk(clk),
    .x(xmulin),
    .r(mulinvlog2_n2729));
  /* fppowbf16.vhdl:4695:44  */
  assign n2733 = {1'b0, absk};
  /* fppowbf16.vhdl:4695:37  */
  assign n2735 = 9'b000000000 - n2733;
  /* fppowbf16.vhdl:4696:19  */
  assign n2736 = xsign_d3 ? minusabsk : n2738;
  /* fppowbf16.vhdl:4696:50  */
  assign n2738 = {1'b0, absk};
  /* fppowbf16.vhdl:4697:4  */
  fixrealkcm_freq500_uid89 mullog2 (
    .clk(clk),
    .x(absk),
    .r(mullog2_n2739));
  /* fppowbf16.vhdl:4701:36  */
  assign n2742 = ufixx[9:0]; // extract
  /* fppowbf16.vhdl:4701:63  */
  assign n2743 = ~xsign_d2;
  /* fppowbf16.vhdl:4701:50  */
  assign n2744 = n2743 ? n2742 : n2746;
  /* fppowbf16.vhdl:4701:100  */
  assign n2745 = ufixx[9:0]; // extract
  /* fppowbf16.vhdl:4701:73  */
  assign n2746 = ~n2745;
  /* fppowbf16.vhdl:4702:22  */
  assign n2747 = absklog2[9:0]; // extract
  /* fppowbf16.vhdl:4702:35  */
  assign n2748 = xsign_d4 ? n2747 : n2750;
  /* fppowbf16.vhdl:4702:71  */
  assign n2749 = absklog2[9:0]; // extract
  /* fppowbf16.vhdl:4702:58  */
  assign n2750 = ~n2749;
  /* fppowbf16.vhdl:4703:4  */
  intadder_10_freq500_uid102 theyadder (
    .clk(clk),
    .x(subop1),
    .y(subop2),
    .cin(n2751),
    .r(theyadder_n2752));
  /* fppowbf16.vhdl:4710:4  */
  fixfunctionbytable_freq500_uid104 expytable (
    .x(y),
    .y(expytable_n2755));
  /* fppowbf16.vhdl:4682:10  */
  always @(posedge clk)
    n2758 <= xsign;
  /* fppowbf16.vhdl:4682:10  */
  always @(posedge clk)
    n2759 <= xsign_d1;
  /* fppowbf16.vhdl:4682:10  */
  always @(posedge clk)
    n2760 <= xsign_d2;
  /* fppowbf16.vhdl:4682:10  */
  always @(posedge clk)
    n2761 <= xsign_d3;
endmodule

module leftshifter19_by_max_16_freq500_uid73
  (input  clk,
   input  [18:0] x,
   input  [4:0] s,
   output [34:0] r);
  wire [4:0] ps;
  wire [4:0] ps_d1;
  wire [18:0] level0;
  wire [18:0] level0_d1;
  wire [19:0] level1;
  wire [21:0] level2;
  wire [25:0] level3;
  wire [25:0] level3_d1;
  wire [33:0] level4;
  wire [49:0] level5;
  wire [19:0] n2685;
  wire n2686;
  wire [19:0] n2687;
  wire [19:0] n2689;
  wire [21:0] n2691;
  wire n2692;
  wire [21:0] n2693;
  wire [21:0] n2695;
  wire [25:0] n2697;
  wire n2698;
  wire [25:0] n2699;
  wire [25:0] n2701;
  wire [33:0] n2703;
  wire n2704;
  wire [33:0] n2705;
  wire [33:0] n2707;
  wire [49:0] n2709;
  wire n2710;
  wire [49:0] n2711;
  wire [49:0] n2713;
  wire [34:0] n2714;
  reg [4:0] n2715;
  reg [18:0] n2716;
  reg [25:0] n2717;
  assign r = n2714; //(module output)
  /* fppowbf16.vhdl:4005:12  */
  assign ps_d1 = n2715; // (signal)
  /* fppowbf16.vhdl:4007:16  */
  assign level0_d1 = n2716; // (signal)
  /* fppowbf16.vhdl:4009:8  */
  assign level1 = n2687; // (signal)
  /* fppowbf16.vhdl:4011:8  */
  assign level2 = n2693; // (signal)
  /* fppowbf16.vhdl:4013:8  */
  assign level3 = n2699; // (signal)
  /* fppowbf16.vhdl:4013:16  */
  assign level3_d1 = n2717; // (signal)
  /* fppowbf16.vhdl:4015:8  */
  assign level4 = n2705; // (signal)
  /* fppowbf16.vhdl:4017:8  */
  assign level5 = n2711; // (signal)
  /* fppowbf16.vhdl:4030:23  */
  assign n2685 = {level0_d1, 1'b0};
  /* fppowbf16.vhdl:4030:52  */
  assign n2686 = ps[0]; // extract
  /* fppowbf16.vhdl:4030:45  */
  assign n2687 = n2686 ? n2685 : n2689;
  /* fppowbf16.vhdl:4030:90  */
  assign n2689 = {1'b0, level0_d1};
  /* fppowbf16.vhdl:4031:20  */
  assign n2691 = {level1, 2'b00};
  /* fppowbf16.vhdl:4031:49  */
  assign n2692 = ps[1]; // extract
  /* fppowbf16.vhdl:4031:42  */
  assign n2693 = n2692 ? n2691 : n2695;
  /* fppowbf16.vhdl:4031:87  */
  assign n2695 = {2'b00, level1};
  /* fppowbf16.vhdl:4032:20  */
  assign n2697 = {level2, 4'b0000};
  /* fppowbf16.vhdl:4032:49  */
  assign n2698 = ps[2]; // extract
  /* fppowbf16.vhdl:4032:42  */
  assign n2699 = n2698 ? n2697 : n2701;
  /* fppowbf16.vhdl:4032:87  */
  assign n2701 = {4'b0000, level2};
  /* fppowbf16.vhdl:4033:23  */
  assign n2703 = {level3_d1, 8'b00000000};
  /* fppowbf16.vhdl:4033:55  */
  assign n2704 = ps_d1[3]; // extract
  /* fppowbf16.vhdl:4033:45  */
  assign n2705 = n2704 ? n2703 : n2707;
  /* fppowbf16.vhdl:4033:93  */
  assign n2707 = {8'b00000000, level3_d1};
  /* fppowbf16.vhdl:4034:20  */
  assign n2709 = {level4, 16'b0000000000000000};
  /* fppowbf16.vhdl:4034:53  */
  assign n2710 = ps_d1[4]; // extract
  /* fppowbf16.vhdl:4034:43  */
  assign n2711 = n2710 ? n2709 : n2713;
  /* fppowbf16.vhdl:4034:92  */
  assign n2713 = {16'b0000000000000000, level4};
  /* fppowbf16.vhdl:4035:15  */
  assign n2714 = level5[34:0]; // extract
  /* fppowbf16.vhdl:4022:10  */
  always @(posedge clk)
    n2715 <= ps;
  /* fppowbf16.vhdl:4022:10  */
  always @(posedge clk)
    n2716 <= level0;
  /* fppowbf16.vhdl:4022:10  */
  always @(posedge clk)
    n2717 <= level3;
endmodule

module intadder_28_freq500_uid69
  (input  clk,
   input  [27:0] x,
   input  [27:0] y,
   input  cin,
   output [27:0] r);
  wire [27:0] rtmp;
  wire [27:0] y_d1;
  wire [27:0] y_d2;
  wire [27:0] y_d3;
  wire [27:0] y_d4;
  wire [27:0] y_d5;
  wire [27:0] y_d6;
  wire [27:0] y_d7;
  wire [27:0] y_d8;
  wire [27:0] y_d9;
  wire [27:0] y_d10;
  wire [27:0] y_d11;
  wire [27:0] y_d12;
  wire [27:0] y_d13;
  wire cin_d1;
  wire cin_d2;
  wire cin_d3;
  wire cin_d4;
  wire cin_d5;
  wire cin_d6;
  wire cin_d7;
  wire cin_d8;
  wire cin_d9;
  wire cin_d10;
  wire cin_d11;
  wire cin_d12;
  wire cin_d13;
  wire [27:0] n2647;
  wire [27:0] n2648;
  wire [27:0] n2649;
  reg [27:0] n2650;
  reg [27:0] n2651;
  reg [27:0] n2652;
  reg [27:0] n2653;
  reg [27:0] n2654;
  reg [27:0] n2655;
  reg [27:0] n2656;
  reg [27:0] n2657;
  reg [27:0] n2658;
  reg [27:0] n2659;
  reg [27:0] n2660;
  reg [27:0] n2661;
  reg [27:0] n2662;
  reg n2663;
  reg n2664;
  reg n2665;
  reg n2666;
  reg n2667;
  reg n2668;
  reg n2669;
  reg n2670;
  reg n2671;
  reg n2672;
  reg n2673;
  reg n2674;
  reg n2675;
  assign r = rtmp; //(module output)
  /* fppowbf16.vhdl:3750:8  */
  assign rtmp = n2649; // (signal)
  /* fppowbf16.vhdl:3752:8  */
  assign y_d1 = n2650; // (signal)
  /* fppowbf16.vhdl:3752:14  */
  assign y_d2 = n2651; // (signal)
  /* fppowbf16.vhdl:3752:20  */
  assign y_d3 = n2652; // (signal)
  /* fppowbf16.vhdl:3752:26  */
  assign y_d4 = n2653; // (signal)
  /* fppowbf16.vhdl:3752:32  */
  assign y_d5 = n2654; // (signal)
  /* fppowbf16.vhdl:3752:38  */
  assign y_d6 = n2655; // (signal)
  /* fppowbf16.vhdl:3752:44  */
  assign y_d7 = n2656; // (signal)
  /* fppowbf16.vhdl:3752:50  */
  assign y_d8 = n2657; // (signal)
  /* fppowbf16.vhdl:3752:56  */
  assign y_d9 = n2658; // (signal)
  /* fppowbf16.vhdl:3752:62  */
  assign y_d10 = n2659; // (signal)
  /* fppowbf16.vhdl:3752:69  */
  assign y_d11 = n2660; // (signal)
  /* fppowbf16.vhdl:3752:76  */
  assign y_d12 = n2661; // (signal)
  /* fppowbf16.vhdl:3752:83  */
  assign y_d13 = n2662; // (signal)
  /* fppowbf16.vhdl:3754:8  */
  assign cin_d1 = n2663; // (signal)
  /* fppowbf16.vhdl:3754:16  */
  assign cin_d2 = n2664; // (signal)
  /* fppowbf16.vhdl:3754:24  */
  assign cin_d3 = n2665; // (signal)
  /* fppowbf16.vhdl:3754:32  */
  assign cin_d4 = n2666; // (signal)
  /* fppowbf16.vhdl:3754:40  */
  assign cin_d5 = n2667; // (signal)
  /* fppowbf16.vhdl:3754:48  */
  assign cin_d6 = n2668; // (signal)
  /* fppowbf16.vhdl:3754:56  */
  assign cin_d7 = n2669; // (signal)
  /* fppowbf16.vhdl:3754:64  */
  assign cin_d8 = n2670; // (signal)
  /* fppowbf16.vhdl:3754:72  */
  assign cin_d9 = n2671; // (signal)
  /* fppowbf16.vhdl:3754:80  */
  assign cin_d10 = n2672; // (signal)
  /* fppowbf16.vhdl:3754:89  */
  assign cin_d11 = n2673; // (signal)
  /* fppowbf16.vhdl:3754:98  */
  assign cin_d12 = n2674; // (signal)
  /* fppowbf16.vhdl:3754:107  */
  assign cin_d13 = n2675; // (signal)
  /* fppowbf16.vhdl:3788:14  */
  assign n2647 = x + y_d13;
  /* fppowbf16.vhdl:3788:22  */
  assign n2648 = {27'b0, cin_d13};  //  uext
  /* fppowbf16.vhdl:3788:22  */
  assign n2649 = n2647 + n2648;
  /* fppowbf16.vhdl:3759:10  */
  always @(posedge clk)
    n2650 <= y;
  /* fppowbf16.vhdl:3759:10  */
  always @(posedge clk)
    n2651 <= y_d1;
  /* fppowbf16.vhdl:3759:10  */
  always @(posedge clk)
    n2652 <= y_d2;
  /* fppowbf16.vhdl:3759:10  */
  always @(posedge clk)
    n2653 <= y_d3;
  /* fppowbf16.vhdl:3759:10  */
  always @(posedge clk)
    n2654 <= y_d4;
  /* fppowbf16.vhdl:3759:10  */
  always @(posedge clk)
    n2655 <= y_d5;
  /* fppowbf16.vhdl:3759:10  */
  always @(posedge clk)
    n2656 <= y_d6;
  /* fppowbf16.vhdl:3759:10  */
  always @(posedge clk)
    n2657 <= y_d7;
  /* fppowbf16.vhdl:3759:10  */
  always @(posedge clk)
    n2658 <= y_d8;
  /* fppowbf16.vhdl:3759:10  */
  always @(posedge clk)
    n2659 <= y_d9;
  /* fppowbf16.vhdl:3759:10  */
  always @(posedge clk)
    n2660 <= y_d10;
  /* fppowbf16.vhdl:3759:10  */
  always @(posedge clk)
    n2661 <= y_d11;
  /* fppowbf16.vhdl:3759:10  */
  always @(posedge clk)
    n2662 <= y_d12;
  /* fppowbf16.vhdl:3759:10  */
  always @(posedge clk)
    n2663 <= cin;
  /* fppowbf16.vhdl:3759:10  */
  always @(posedge clk)
    n2664 <= cin_d1;
  /* fppowbf16.vhdl:3759:10  */
  always @(posedge clk)
    n2665 <= cin_d2;
  /* fppowbf16.vhdl:3759:10  */
  always @(posedge clk)
    n2666 <= cin_d3;
  /* fppowbf16.vhdl:3759:10  */
  always @(posedge clk)
    n2667 <= cin_d4;
  /* fppowbf16.vhdl:3759:10  */
  always @(posedge clk)
    n2668 <= cin_d5;
  /* fppowbf16.vhdl:3759:10  */
  always @(posedge clk)
    n2669 <= cin_d6;
  /* fppowbf16.vhdl:3759:10  */
  always @(posedge clk)
    n2670 <= cin_d7;
  /* fppowbf16.vhdl:3759:10  */
  always @(posedge clk)
    n2671 <= cin_d8;
  /* fppowbf16.vhdl:3759:10  */
  always @(posedge clk)
    n2672 <= cin_d9;
  /* fppowbf16.vhdl:3759:10  */
  always @(posedge clk)
    n2673 <= cin_d10;
  /* fppowbf16.vhdl:3759:10  */
  always @(posedge clk)
    n2674 <= cin_d11;
  /* fppowbf16.vhdl:3759:10  */
  always @(posedge clk)
    n2675 <= cin_d12;
endmodule

module intmultiplier_18x8_21_freq500_uid65
  (input  clk,
   input  [17:0] x,
   input  [7:0] y,
   output [20:0] r);
  wire [17:0] xx;
  wire [7:0] yy;
  wire [7:0] yy_d1;
  wire [7:0] yy_d2;
  wire [7:0] yy_d3;
  wire [7:0] yy_d4;
  wire [7:0] yy_d5;
  wire [7:0] yy_d6;
  wire [7:0] yy_d7;
  wire [7:0] yy_d8;
  wire [7:0] yy_d9;
  wire [7:0] yy_d10;
  wire [7:0] yy_d11;
  wire [25:0] rr;
  wire [25:0] n2601;
  wire [25:0] n2602;
  wire [25:0] n2603;
  wire [20:0] n2604;
  reg [7:0] n2605;
  reg [7:0] n2606;
  reg [7:0] n2607;
  reg [7:0] n2608;
  reg [7:0] n2609;
  reg [7:0] n2610;
  reg [7:0] n2611;
  reg [7:0] n2612;
  reg [7:0] n2613;
  reg [7:0] n2614;
  reg [7:0] n2615;
  assign r = n2604; //(module output)
  /* fppowbf16.vhdl:3689:12  */
  assign yy_d1 = n2605; // (signal)
  /* fppowbf16.vhdl:3689:19  */
  assign yy_d2 = n2606; // (signal)
  /* fppowbf16.vhdl:3689:26  */
  assign yy_d3 = n2607; // (signal)
  /* fppowbf16.vhdl:3689:33  */
  assign yy_d4 = n2608; // (signal)
  /* fppowbf16.vhdl:3689:40  */
  assign yy_d5 = n2609; // (signal)
  /* fppowbf16.vhdl:3689:47  */
  assign yy_d6 = n2610; // (signal)
  /* fppowbf16.vhdl:3689:54  */
  assign yy_d7 = n2611; // (signal)
  /* fppowbf16.vhdl:3689:61  */
  assign yy_d8 = n2612; // (signal)
  /* fppowbf16.vhdl:3689:68  */
  assign yy_d9 = n2613; // (signal)
  /* fppowbf16.vhdl:3689:75  */
  assign yy_d10 = n2614; // (signal)
  /* fppowbf16.vhdl:3689:83  */
  assign yy_d11 = n2615; // (signal)
  /* fppowbf16.vhdl:3691:8  */
  assign rr = n2603; // (signal)
  /* fppowbf16.vhdl:3714:12  */
  assign n2601 = {8'b0, xx};  //  uext
  /* fppowbf16.vhdl:3714:12  */
  assign n2602 = {18'b0, yy_d11};  //  uext
  /* fppowbf16.vhdl:3714:12  */
  assign n2603 = n2601 * n2602; // umul
  /* fppowbf16.vhdl:3715:28  */
  assign n2604 = rr[25:5]; // extract
  /* fppowbf16.vhdl:3696:10  */
  always @(posedge clk)
    n2605 <= yy;
  /* fppowbf16.vhdl:3696:10  */
  always @(posedge clk)
    n2606 <= yy_d1;
  /* fppowbf16.vhdl:3696:10  */
  always @(posedge clk)
    n2607 <= yy_d2;
  /* fppowbf16.vhdl:3696:10  */
  always @(posedge clk)
    n2608 <= yy_d3;
  /* fppowbf16.vhdl:3696:10  */
  always @(posedge clk)
    n2609 <= yy_d4;
  /* fppowbf16.vhdl:3696:10  */
  always @(posedge clk)
    n2610 <= yy_d5;
  /* fppowbf16.vhdl:3696:10  */
  always @(posedge clk)
    n2611 <= yy_d6;
  /* fppowbf16.vhdl:3696:10  */
  always @(posedge clk)
    n2612 <= yy_d7;
  /* fppowbf16.vhdl:3696:10  */
  always @(posedge clk)
    n2613 <= yy_d8;
  /* fppowbf16.vhdl:3696:10  */
  always @(posedge clk)
    n2614 <= yy_d9;
  /* fppowbf16.vhdl:3696:10  */
  always @(posedge clk)
    n2615 <= yy_d10;
endmodule

module intadder_25_freq500_uid60
  (input  clk,
   input  [24:0] x,
   input  [24:0] y,
   input  cin,
   output [24:0] r);
  wire [24:0] rtmp;
  wire cin_d1;
  wire cin_d2;
  wire cin_d3;
  wire cin_d4;
  wire cin_d5;
  wire cin_d6;
  wire cin_d7;
  wire cin_d8;
  wire cin_d9;
  wire cin_d10;
  wire cin_d11;
  wire [24:0] n2571;
  wire [24:0] n2572;
  wire [24:0] n2573;
  reg n2574;
  reg n2575;
  reg n2576;
  reg n2577;
  reg n2578;
  reg n2579;
  reg n2580;
  reg n2581;
  reg n2582;
  reg n2583;
  reg n2584;
  assign r = rtmp; //(module output)
  /* fppowbf16.vhdl:3066:8  */
  assign rtmp = n2573; // (signal)
  /* fppowbf16.vhdl:3068:8  */
  assign cin_d1 = n2574; // (signal)
  /* fppowbf16.vhdl:3068:16  */
  assign cin_d2 = n2575; // (signal)
  /* fppowbf16.vhdl:3068:24  */
  assign cin_d3 = n2576; // (signal)
  /* fppowbf16.vhdl:3068:32  */
  assign cin_d4 = n2577; // (signal)
  /* fppowbf16.vhdl:3068:40  */
  assign cin_d5 = n2578; // (signal)
  /* fppowbf16.vhdl:3068:48  */
  assign cin_d6 = n2579; // (signal)
  /* fppowbf16.vhdl:3068:56  */
  assign cin_d7 = n2580; // (signal)
  /* fppowbf16.vhdl:3068:64  */
  assign cin_d8 = n2581; // (signal)
  /* fppowbf16.vhdl:3068:72  */
  assign cin_d9 = n2582; // (signal)
  /* fppowbf16.vhdl:3068:80  */
  assign cin_d10 = n2583; // (signal)
  /* fppowbf16.vhdl:3068:89  */
  assign cin_d11 = n2584; // (signal)
  /* fppowbf16.vhdl:3087:14  */
  assign n2571 = x + y;
  /* fppowbf16.vhdl:3087:18  */
  assign n2572 = {24'b0, cin_d11};  //  uext
  /* fppowbf16.vhdl:3087:18  */
  assign n2573 = n2571 + n2572;
  /* fppowbf16.vhdl:3073:10  */
  always @(posedge clk)
    n2574 <= cin;
  /* fppowbf16.vhdl:3073:10  */
  always @(posedge clk)
    n2575 <= cin_d1;
  /* fppowbf16.vhdl:3073:10  */
  always @(posedge clk)
    n2576 <= cin_d2;
  /* fppowbf16.vhdl:3073:10  */
  always @(posedge clk)
    n2577 <= cin_d3;
  /* fppowbf16.vhdl:3073:10  */
  always @(posedge clk)
    n2578 <= cin_d4;
  /* fppowbf16.vhdl:3073:10  */
  always @(posedge clk)
    n2579 <= cin_d5;
  /* fppowbf16.vhdl:3073:10  */
  always @(posedge clk)
    n2580 <= cin_d6;
  /* fppowbf16.vhdl:3073:10  */
  always @(posedge clk)
    n2581 <= cin_d7;
  /* fppowbf16.vhdl:3073:10  */
  always @(posedge clk)
    n2582 <= cin_d8;
  /* fppowbf16.vhdl:3073:10  */
  always @(posedge clk)
    n2583 <= cin_d9;
  /* fppowbf16.vhdl:3073:10  */
  always @(posedge clk)
    n2584 <= cin_d10;
endmodule

module intadder_23_freq500_uid57
  (input  clk,
   input  [22:0] x,
   input  [22:0] y,
   input  cin,
   output [22:0] r);
  wire [22:0] rtmp;
  wire [22:0] x_d1;
  wire [22:0] x_d2;
  wire cin_d1;
  wire cin_d2;
  wire cin_d3;
  wire cin_d4;
  wire cin_d5;
  wire cin_d6;
  wire [22:0] n2544;
  wire [22:0] n2545;
  wire [22:0] n2546;
  reg [22:0] n2547;
  reg [22:0] n2548;
  reg n2549;
  reg n2550;
  reg n2551;
  reg n2552;
  reg n2553;
  reg n2554;
  assign r = rtmp; //(module output)
  /* fppowbf16.vhdl:3010:8  */
  assign rtmp = n2546; // (signal)
  /* fppowbf16.vhdl:3012:8  */
  assign x_d1 = n2547; // (signal)
  /* fppowbf16.vhdl:3012:14  */
  assign x_d2 = n2548; // (signal)
  /* fppowbf16.vhdl:3014:8  */
  assign cin_d1 = n2549; // (signal)
  /* fppowbf16.vhdl:3014:16  */
  assign cin_d2 = n2550; // (signal)
  /* fppowbf16.vhdl:3014:24  */
  assign cin_d3 = n2551; // (signal)
  /* fppowbf16.vhdl:3014:32  */
  assign cin_d4 = n2552; // (signal)
  /* fppowbf16.vhdl:3014:40  */
  assign cin_d5 = n2553; // (signal)
  /* fppowbf16.vhdl:3014:48  */
  assign cin_d6 = n2554; // (signal)
  /* fppowbf16.vhdl:3030:17  */
  assign n2544 = x_d2 + y;
  /* fppowbf16.vhdl:3030:21  */
  assign n2545 = {22'b0, cin_d6};  //  uext
  /* fppowbf16.vhdl:3030:21  */
  assign n2546 = n2544 + n2545;
  /* fppowbf16.vhdl:3019:10  */
  always @(posedge clk)
    n2547 <= x;
  /* fppowbf16.vhdl:3019:10  */
  always @(posedge clk)
    n2548 <= x_d1;
  /* fppowbf16.vhdl:3019:10  */
  always @(posedge clk)
    n2549 <= cin;
  /* fppowbf16.vhdl:3019:10  */
  always @(posedge clk)
    n2550 <= cin_d1;
  /* fppowbf16.vhdl:3019:10  */
  always @(posedge clk)
    n2551 <= cin_d2;
  /* fppowbf16.vhdl:3019:10  */
  always @(posedge clk)
    n2552 <= cin_d3;
  /* fppowbf16.vhdl:3019:10  */
  always @(posedge clk)
    n2553 <= cin_d4;
  /* fppowbf16.vhdl:3019:10  */
  always @(posedge clk)
    n2554 <= cin_d5;
endmodule

module rightshifter14_by_max_13_freq500_uid55
  (input  clk,
   input  [13:0] x,
   input  [3:0] s,
   output [26:0] r);
  wire [3:0] ps;
  wire [3:0] ps_d1;
  wire [3:0] ps_d2;
  wire [3:0] ps_d3;
  wire [13:0] level0;
  wire [14:0] level1;
  wire [16:0] level2;
  wire [20:0] level3;
  wire [20:0] level3_d1;
  wire [28:0] level4;
  wire [14:0] n2503;
  wire n2504;
  wire [14:0] n2505;
  wire [14:0] n2507;
  wire [16:0] n2509;
  wire n2510;
  wire [16:0] n2511;
  wire [16:0] n2513;
  wire [20:0] n2515;
  wire n2516;
  wire [20:0] n2517;
  wire [20:0] n2519;
  wire [28:0] n2521;
  wire n2522;
  wire [28:0] n2523;
  wire [28:0] n2525;
  wire [26:0] n2526;
  reg [3:0] n2527;
  reg [3:0] n2528;
  reg [3:0] n2529;
  reg [20:0] n2530;
  assign r = n2526; //(module output)
  /* fppowbf16.vhdl:2947:12  */
  assign ps_d1 = n2527; // (signal)
  /* fppowbf16.vhdl:2947:19  */
  assign ps_d2 = n2528; // (signal)
  /* fppowbf16.vhdl:2947:26  */
  assign ps_d3 = n2529; // (signal)
  /* fppowbf16.vhdl:2951:8  */
  assign level1 = n2505; // (signal)
  /* fppowbf16.vhdl:2953:8  */
  assign level2 = n2511; // (signal)
  /* fppowbf16.vhdl:2955:8  */
  assign level3 = n2517; // (signal)
  /* fppowbf16.vhdl:2955:16  */
  assign level3_d1 = n2530; // (signal)
  /* fppowbf16.vhdl:2957:8  */
  assign level4 = n2523; // (signal)
  /* fppowbf16.vhdl:2971:35  */
  assign n2503 = {1'b0, level0};
  /* fppowbf16.vhdl:2971:54  */
  assign n2504 = ps_d2[0]; // extract
  /* fppowbf16.vhdl:2971:44  */
  assign n2505 = n2504 ? n2503 : n2507;
  /* fppowbf16.vhdl:2971:79  */
  assign n2507 = {level0, 1'b0};
  /* fppowbf16.vhdl:2972:35  */
  assign n2509 = {2'b00, level1};
  /* fppowbf16.vhdl:2972:54  */
  assign n2510 = ps_d2[1]; // extract
  /* fppowbf16.vhdl:2972:44  */
  assign n2511 = n2510 ? n2509 : n2513;
  /* fppowbf16.vhdl:2972:79  */
  assign n2513 = {level1, 2'b00};
  /* fppowbf16.vhdl:2973:35  */
  assign n2515 = {4'b0000, level2};
  /* fppowbf16.vhdl:2973:54  */
  assign n2516 = ps_d2[2]; // extract
  /* fppowbf16.vhdl:2973:44  */
  assign n2517 = n2516 ? n2515 : n2519;
  /* fppowbf16.vhdl:2973:79  */
  assign n2519 = {level2, 4'b0000};
  /* fppowbf16.vhdl:2974:35  */
  assign n2521 = {8'b00000000, level3_d1};
  /* fppowbf16.vhdl:2974:57  */
  assign n2522 = ps_d3[3]; // extract
  /* fppowbf16.vhdl:2974:47  */
  assign n2523 = n2522 ? n2521 : n2525;
  /* fppowbf16.vhdl:2974:85  */
  assign n2525 = {level3_d1, 8'b00000000};
  /* fppowbf16.vhdl:2975:15  */
  assign n2526 = level4[28:2]; // extract
  /* fppowbf16.vhdl:2962:10  */
  always @(posedge clk)
    n2527 <= ps;
  /* fppowbf16.vhdl:2962:10  */
  always @(posedge clk)
    n2528 <= ps_d1;
  /* fppowbf16.vhdl:2962:10  */
  always @(posedge clk)
    n2529 <= ps_d2;
  /* fppowbf16.vhdl:2962:10  */
  always @(posedge clk)
    n2530 <= level3;
endmodule

module normalizer_z_38_30_16_freq500_uid53
  (input  clk,
   input  [37:0] x,
   output [4:0] count,
   output [29:0] r);
  wire [37:0] level5;
  wire count4;
  wire count4_d1;
  wire count4_d2;
  wire [37:0] level4;
  wire [37:0] level4_d1;
  wire count3;
  wire count3_d1;
  wire [36:0] level3;
  wire count2;
  wire count2_d1;
  wire [32:0] level2;
  wire [32:0] level2_d1;
  wire count1;
  wire [30:0] level1;
  wire [30:0] level1_d1;
  wire count0;
  wire count0_d1;
  wire [29:0] level0;
  wire [4:0] scount;
  wire [15:0] n2429;
  wire n2431;
  wire n2432;
  wire n2434;
  wire [37:0] n2435;
  wire [21:0] n2436;
  wire [37:0] n2438;
  wire [7:0] n2440;
  wire n2442;
  wire n2443;
  wire [36:0] n2445;
  wire n2446;
  wire [36:0] n2447;
  wire [29:0] n2448;
  wire [36:0] n2450;
  wire [3:0] n2452;
  wire n2454;
  wire n2455;
  wire [32:0] n2457;
  wire n2458;
  wire [32:0] n2459;
  wire [32:0] n2460;
  wire [1:0] n2462;
  wire n2464;
  wire n2465;
  wire [30:0] n2467;
  wire n2468;
  wire [30:0] n2469;
  wire [30:0] n2470;
  wire n2472;
  wire n2474;
  wire n2475;
  wire [29:0] n2477;
  wire n2478;
  wire [29:0] n2479;
  wire [29:0] n2480;
  wire [1:0] n2481;
  wire [2:0] n2482;
  wire [3:0] n2483;
  wire [4:0] n2484;
  reg n2485;
  reg n2486;
  reg [37:0] n2487;
  reg n2488;
  reg n2489;
  reg [32:0] n2490;
  reg [30:0] n2491;
  reg n2492;
  assign count = scount; //(module output)
  assign r = level0; //(module output)
  /* fppowbf16.vhdl:2859:8  */
  assign count4 = n2432; // (signal)
  /* fppowbf16.vhdl:2859:16  */
  assign count4_d1 = n2485; // (signal)
  /* fppowbf16.vhdl:2859:27  */
  assign count4_d2 = n2486; // (signal)
  /* fppowbf16.vhdl:2861:8  */
  assign level4 = n2435; // (signal)
  /* fppowbf16.vhdl:2861:16  */
  assign level4_d1 = n2487; // (signal)
  /* fppowbf16.vhdl:2863:8  */
  assign count3 = n2443; // (signal)
  /* fppowbf16.vhdl:2863:16  */
  assign count3_d1 = n2488; // (signal)
  /* fppowbf16.vhdl:2865:8  */
  assign level3 = n2447; // (signal)
  /* fppowbf16.vhdl:2867:8  */
  assign count2 = n2455; // (signal)
  /* fppowbf16.vhdl:2867:16  */
  assign count2_d1 = n2489; // (signal)
  /* fppowbf16.vhdl:2869:8  */
  assign level2 = n2459; // (signal)
  /* fppowbf16.vhdl:2869:16  */
  assign level2_d1 = n2490; // (signal)
  /* fppowbf16.vhdl:2871:8  */
  assign count1 = n2465; // (signal)
  /* fppowbf16.vhdl:2873:8  */
  assign level1 = n2469; // (signal)
  /* fppowbf16.vhdl:2873:16  */
  assign level1_d1 = n2491; // (signal)
  /* fppowbf16.vhdl:2875:8  */
  assign count0 = n2475; // (signal)
  /* fppowbf16.vhdl:2875:16  */
  assign count0_d1 = n2492; // (signal)
  /* fppowbf16.vhdl:2877:8  */
  assign level0 = n2479; // (signal)
  /* fppowbf16.vhdl:2879:8  */
  assign scount = n2484; // (signal)
  /* fppowbf16.vhdl:2896:28  */
  assign n2429 = level5[37:22]; // extract
  /* fppowbf16.vhdl:2896:43  */
  assign n2431 = n2429 == 16'b0000000000000000;
  /* fppowbf16.vhdl:2896:17  */
  assign n2432 = n2431 ? 1'b1 : 1'b0;
  /* fppowbf16.vhdl:2897:44  */
  assign n2434 = ~count4;
  /* fppowbf16.vhdl:2897:33  */
  assign n2435 = n2434 ? level5 : n2438;
  /* fppowbf16.vhdl:2897:60  */
  assign n2436 = level5[21:0]; // extract
  /* fppowbf16.vhdl:2897:74  */
  assign n2438 = {n2436, 16'b0000000000000000};
  /* fppowbf16.vhdl:2899:31  */
  assign n2440 = level4_d1[37:30]; // extract
  /* fppowbf16.vhdl:2899:46  */
  assign n2442 = n2440 == 8'b00000000;
  /* fppowbf16.vhdl:2899:17  */
  assign n2443 = n2442 ? 1'b1 : 1'b0;
  /* fppowbf16.vhdl:2900:22  */
  assign n2445 = level4_d1[37:1]; // extract
  /* fppowbf16.vhdl:2900:47  */
  assign n2446 = ~count3;
  /* fppowbf16.vhdl:2900:36  */
  assign n2447 = n2446 ? n2445 : n2450;
  /* fppowbf16.vhdl:2900:66  */
  assign n2448 = level4_d1[29:0]; // extract
  /* fppowbf16.vhdl:2900:80  */
  assign n2450 = {n2448, 7'b0000000};
  /* fppowbf16.vhdl:2902:28  */
  assign n2452 = level3[36:33]; // extract
  /* fppowbf16.vhdl:2902:43  */
  assign n2454 = n2452 == 4'b0000;
  /* fppowbf16.vhdl:2902:17  */
  assign n2455 = n2454 ? 1'b1 : 1'b0;
  /* fppowbf16.vhdl:2903:19  */
  assign n2457 = level3[36:4]; // extract
  /* fppowbf16.vhdl:2903:44  */
  assign n2458 = ~count2;
  /* fppowbf16.vhdl:2903:33  */
  assign n2459 = n2458 ? n2457 : n2460;
  /* fppowbf16.vhdl:2903:60  */
  assign n2460 = level3[32:0]; // extract
  /* fppowbf16.vhdl:2905:31  */
  assign n2462 = level2_d1[32:31]; // extract
  /* fppowbf16.vhdl:2905:46  */
  assign n2464 = n2462 == 2'b00;
  /* fppowbf16.vhdl:2905:17  */
  assign n2465 = n2464 ? 1'b1 : 1'b0;
  /* fppowbf16.vhdl:2906:22  */
  assign n2467 = level2_d1[32:2]; // extract
  /* fppowbf16.vhdl:2906:47  */
  assign n2468 = ~count1;
  /* fppowbf16.vhdl:2906:36  */
  assign n2469 = n2468 ? n2467 : n2470;
  /* fppowbf16.vhdl:2906:66  */
  assign n2470 = level2_d1[30:0]; // extract
  /* fppowbf16.vhdl:2908:28  */
  assign n2472 = level1[30]; // extract
  /* fppowbf16.vhdl:2908:43  */
  assign n2474 = n2472 == 1'b0;
  /* fppowbf16.vhdl:2908:17  */
  assign n2475 = n2474 ? 1'b1 : 1'b0;
  /* fppowbf16.vhdl:2909:22  */
  assign n2477 = level1_d1[30:1]; // extract
  /* fppowbf16.vhdl:2909:50  */
  assign n2478 = ~count0_d1;
  /* fppowbf16.vhdl:2909:36  */
  assign n2479 = n2478 ? n2477 : n2480;
  /* fppowbf16.vhdl:2909:69  */
  assign n2480 = level1_d1[29:0]; // extract
  /* fppowbf16.vhdl:2912:24  */
  assign n2481 = {count4_d2, count3_d1};
  /* fppowbf16.vhdl:2912:36  */
  assign n2482 = {n2481, count2_d1};
  /* fppowbf16.vhdl:2912:48  */
  assign n2483 = {n2482, count1};
  /* fppowbf16.vhdl:2912:57  */
  assign n2484 = {n2483, count0};
  /* fppowbf16.vhdl:2884:10  */
  always @(posedge clk)
    n2485 <= count4;
  /* fppowbf16.vhdl:2884:10  */
  always @(posedge clk)
    n2486 <= count4_d1;
  /* fppowbf16.vhdl:2884:10  */
  always @(posedge clk)
    n2487 <= level4;
  /* fppowbf16.vhdl:2884:10  */
  always @(posedge clk)
    n2488 <= count3;
  /* fppowbf16.vhdl:2884:10  */
  always @(posedge clk)
    n2489 <= count2;
  /* fppowbf16.vhdl:2884:10  */
  always @(posedge clk)
    n2490 <= level2;
  /* fppowbf16.vhdl:2884:10  */
  always @(posedge clk)
    n2491 <= level1;
  /* fppowbf16.vhdl:2884:10  */
  always @(posedge clk)
    n2492 <= count0;
endmodule

module intadder_38_freq500_uid51
  (input  clk,
   input  [37:0] x,
   input  [37:0] y,
   input  cin,
   output [37:0] r);
  wire cin_0;
  wire cin_0_d1;
  wire cin_0_d2;
  wire cin_0_d3;
  wire cin_0_d4;
  wire cin_0_d5;
  wire cin_0_d6;
  wire cin_0_d7;
  wire [25:0] x_0;
  wire [25:0] x_0_d1;
  wire [25:0] x_0_d2;
  wire [25:0] x_0_d3;
  wire [25:0] x_0_d4;
  wire [25:0] x_0_d5;
  wire [25:0] x_0_d6;
  wire [25:0] y_0;
  wire [25:0] y_0_d1;
  wire [25:0] s_0;
  wire [24:0] r_0;
  wire [24:0] r_0_d1;
  wire cin_1;
  wire cin_1_d1;
  wire [13:0] x_1;
  wire [13:0] x_1_d1;
  wire [13:0] x_1_d2;
  wire [13:0] x_1_d3;
  wire [13:0] x_1_d4;
  wire [13:0] x_1_d5;
  wire [13:0] x_1_d6;
  wire [13:0] x_1_d7;
  wire [13:0] y_1;
  wire [13:0] y_1_d1;
  wire [13:0] y_1_d2;
  wire [13:0] s_1;
  wire [12:0] r_1;
  wire [24:0] n2367;
  wire [25:0] n2369;
  wire [24:0] n2370;
  wire [25:0] n2372;
  wire [25:0] n2373;
  wire [25:0] n2374;
  wire [25:0] n2375;
  wire [24:0] n2376;
  wire n2377;
  wire [12:0] n2378;
  wire [13:0] n2380;
  wire [12:0] n2381;
  wire [13:0] n2383;
  wire [13:0] n2384;
  wire [13:0] n2385;
  wire [13:0] n2386;
  wire [12:0] n2387;
  wire [37:0] n2388;
  reg n2389;
  reg n2390;
  reg n2391;
  reg n2392;
  reg n2393;
  reg n2394;
  reg n2395;
  reg [25:0] n2396;
  reg [25:0] n2397;
  reg [25:0] n2398;
  reg [25:0] n2399;
  reg [25:0] n2400;
  reg [25:0] n2401;
  reg [25:0] n2402;
  reg [24:0] n2403;
  reg n2404;
  reg [13:0] n2405;
  reg [13:0] n2406;
  reg [13:0] n2407;
  reg [13:0] n2408;
  reg [13:0] n2409;
  reg [13:0] n2410;
  reg [13:0] n2411;
  reg [13:0] n2412;
  reg [13:0] n2413;
  assign r = n2388; //(module output)
  /* fppowbf16.vhdl:2762:15  */
  assign cin_0_d1 = n2389; // (signal)
  /* fppowbf16.vhdl:2762:25  */
  assign cin_0_d2 = n2390; // (signal)
  /* fppowbf16.vhdl:2762:35  */
  assign cin_0_d3 = n2391; // (signal)
  /* fppowbf16.vhdl:2762:45  */
  assign cin_0_d4 = n2392; // (signal)
  /* fppowbf16.vhdl:2762:55  */
  assign cin_0_d5 = n2393; // (signal)
  /* fppowbf16.vhdl:2762:65  */
  assign cin_0_d6 = n2394; // (signal)
  /* fppowbf16.vhdl:2762:75  */
  assign cin_0_d7 = n2395; // (signal)
  /* fppowbf16.vhdl:2764:8  */
  assign x_0 = n2369; // (signal)
  /* fppowbf16.vhdl:2764:13  */
  assign x_0_d1 = n2396; // (signal)
  /* fppowbf16.vhdl:2764:21  */
  assign x_0_d2 = n2397; // (signal)
  /* fppowbf16.vhdl:2764:29  */
  assign x_0_d3 = n2398; // (signal)
  /* fppowbf16.vhdl:2764:37  */
  assign x_0_d4 = n2399; // (signal)
  /* fppowbf16.vhdl:2764:45  */
  assign x_0_d5 = n2400; // (signal)
  /* fppowbf16.vhdl:2764:53  */
  assign x_0_d6 = n2401; // (signal)
  /* fppowbf16.vhdl:2766:8  */
  assign y_0 = n2372; // (signal)
  /* fppowbf16.vhdl:2766:13  */
  assign y_0_d1 = n2402; // (signal)
  /* fppowbf16.vhdl:2768:8  */
  assign s_0 = n2375; // (signal)
  /* fppowbf16.vhdl:2770:8  */
  assign r_0 = n2376; // (signal)
  /* fppowbf16.vhdl:2770:13  */
  assign r_0_d1 = n2403; // (signal)
  /* fppowbf16.vhdl:2772:8  */
  assign cin_1 = n2377; // (signal)
  /* fppowbf16.vhdl:2772:15  */
  assign cin_1_d1 = n2404; // (signal)
  /* fppowbf16.vhdl:2774:8  */
  assign x_1 = n2380; // (signal)
  /* fppowbf16.vhdl:2774:13  */
  assign x_1_d1 = n2405; // (signal)
  /* fppowbf16.vhdl:2774:21  */
  assign x_1_d2 = n2406; // (signal)
  /* fppowbf16.vhdl:2774:29  */
  assign x_1_d3 = n2407; // (signal)
  /* fppowbf16.vhdl:2774:37  */
  assign x_1_d4 = n2408; // (signal)
  /* fppowbf16.vhdl:2774:45  */
  assign x_1_d5 = n2409; // (signal)
  /* fppowbf16.vhdl:2774:53  */
  assign x_1_d6 = n2410; // (signal)
  /* fppowbf16.vhdl:2774:61  */
  assign x_1_d7 = n2411; // (signal)
  /* fppowbf16.vhdl:2776:8  */
  assign y_1 = n2383; // (signal)
  /* fppowbf16.vhdl:2776:13  */
  assign y_1_d1 = n2412; // (signal)
  /* fppowbf16.vhdl:2776:21  */
  assign y_1_d2 = n2413; // (signal)
  /* fppowbf16.vhdl:2778:8  */
  assign s_1 = n2386; // (signal)
  /* fppowbf16.vhdl:2780:8  */
  assign r_1 = n2387; // (signal)
  /* fppowbf16.vhdl:2814:18  */
  assign n2367 = x[24:0]; // extract
  /* fppowbf16.vhdl:2814:15  */
  assign n2369 = {1'b0, n2367};
  /* fppowbf16.vhdl:2815:18  */
  assign n2370 = y[24:0]; // extract
  /* fppowbf16.vhdl:2815:15  */
  assign n2372 = {1'b0, n2370};
  /* fppowbf16.vhdl:2816:18  */
  assign n2373 = x_0_d6 + y_0_d1;
  /* fppowbf16.vhdl:2816:27  */
  assign n2374 = {25'b0, cin_0_d7};  //  uext
  /* fppowbf16.vhdl:2816:27  */
  assign n2375 = n2373 + n2374;
  /* fppowbf16.vhdl:2817:14  */
  assign n2376 = s_0[24:0]; // extract
  /* fppowbf16.vhdl:2818:16  */
  assign n2377 = s_0[25]; // extract
  /* fppowbf16.vhdl:2819:18  */
  assign n2378 = x[37:25]; // extract
  /* fppowbf16.vhdl:2819:15  */
  assign n2380 = {1'b0, n2378};
  /* fppowbf16.vhdl:2820:18  */
  assign n2381 = y[37:25]; // extract
  /* fppowbf16.vhdl:2820:15  */
  assign n2383 = {1'b0, n2381};
  /* fppowbf16.vhdl:2821:18  */
  assign n2384 = x_1_d7 + y_1_d2;
  /* fppowbf16.vhdl:2821:27  */
  assign n2385 = {13'b0, cin_1_d1};  //  uext
  /* fppowbf16.vhdl:2821:27  */
  assign n2386 = n2384 + n2385;
  /* fppowbf16.vhdl:2822:14  */
  assign n2387 = s_1[12:0]; // extract
  /* fppowbf16.vhdl:2823:13  */
  assign n2388 = {r_1, r_0_d1};
  /* fppowbf16.vhdl:2785:10  */
  always @(posedge clk)
    n2389 <= cin_0;
  /* fppowbf16.vhdl:2785:10  */
  always @(posedge clk)
    n2390 <= cin_0_d1;
  /* fppowbf16.vhdl:2785:10  */
  always @(posedge clk)
    n2391 <= cin_0_d2;
  /* fppowbf16.vhdl:2785:10  */
  always @(posedge clk)
    n2392 <= cin_0_d3;
  /* fppowbf16.vhdl:2785:10  */
  always @(posedge clk)
    n2393 <= cin_0_d4;
  /* fppowbf16.vhdl:2785:10  */
  always @(posedge clk)
    n2394 <= cin_0_d5;
  /* fppowbf16.vhdl:2785:10  */
  always @(posedge clk)
    n2395 <= cin_0_d6;
  /* fppowbf16.vhdl:2785:10  */
  always @(posedge clk)
    n2396 <= x_0;
  /* fppowbf16.vhdl:2785:10  */
  always @(posedge clk)
    n2397 <= x_0_d1;
  /* fppowbf16.vhdl:2785:10  */
  always @(posedge clk)
    n2398 <= x_0_d2;
  /* fppowbf16.vhdl:2785:10  */
  always @(posedge clk)
    n2399 <= x_0_d3;
  /* fppowbf16.vhdl:2785:10  */
  always @(posedge clk)
    n2400 <= x_0_d4;
  /* fppowbf16.vhdl:2785:10  */
  always @(posedge clk)
    n2401 <= x_0_d5;
  /* fppowbf16.vhdl:2785:10  */
  always @(posedge clk)
    n2402 <= y_0;
  /* fppowbf16.vhdl:2785:10  */
  always @(posedge clk)
    n2403 <= r_0;
  /* fppowbf16.vhdl:2785:10  */
  always @(posedge clk)
    n2404 <= cin_1;
  /* fppowbf16.vhdl:2785:10  */
  always @(posedge clk)
    n2405 <= x_1;
  /* fppowbf16.vhdl:2785:10  */
  always @(posedge clk)
    n2406 <= x_1_d1;
  /* fppowbf16.vhdl:2785:10  */
  always @(posedge clk)
    n2407 <= x_1_d2;
  /* fppowbf16.vhdl:2785:10  */
  always @(posedge clk)
    n2408 <= x_1_d3;
  /* fppowbf16.vhdl:2785:10  */
  always @(posedge clk)
    n2409 <= x_1_d4;
  /* fppowbf16.vhdl:2785:10  */
  always @(posedge clk)
    n2410 <= x_1_d5;
  /* fppowbf16.vhdl:2785:10  */
  always @(posedge clk)
    n2411 <= x_1_d6;
  /* fppowbf16.vhdl:2785:10  */
  always @(posedge clk)
    n2412 <= y_1;
  /* fppowbf16.vhdl:2785:10  */
  always @(posedge clk)
    n2413 <= y_1_d1;
endmodule

module fixrealkcm_freq500_uid39
  (input  clk,
   input  [7:0] x,
   output [28:0] r);
  wire [4:0] fixrealkcm_freq500_uid39_a0;
  wire [28:0] fixrealkcm_freq500_uid39_t0;
  wire [28:0] fixrealkcm_freq500_uid39_t0_copy43;
  wire [28:0] fixrealkcm_freq500_uid39_t0_copy43_d1;
  wire bh40_w0_0;
  wire bh40_w1_0;
  wire bh40_w2_0;
  wire bh40_w3_0;
  wire bh40_w4_0;
  wire bh40_w5_0;
  wire bh40_w6_0;
  wire bh40_w7_0;
  wire bh40_w8_0;
  wire bh40_w9_0;
  wire bh40_w10_0;
  wire bh40_w11_0;
  wire bh40_w12_0;
  wire bh40_w13_0;
  wire bh40_w14_0;
  wire bh40_w15_0;
  wire bh40_w16_0;
  wire bh40_w17_0;
  wire bh40_w18_0;
  wire bh40_w19_0;
  wire bh40_w20_0;
  wire bh40_w21_0;
  wire bh40_w22_0;
  wire bh40_w23_0;
  wire bh40_w24_0;
  wire bh40_w25_0;
  wire bh40_w26_0;
  wire bh40_w27_0;
  wire bh40_w28_0;
  wire [2:0] fixrealkcm_freq500_uid39_a1;
  wire [23:0] fixrealkcm_freq500_uid39_t1;
  wire [23:0] fixrealkcm_freq500_uid39_t1_copy46;
  wire [23:0] fixrealkcm_freq500_uid39_t1_copy46_d1;
  wire bh40_w0_1;
  wire bh40_w1_1;
  wire bh40_w2_1;
  wire bh40_w3_1;
  wire bh40_w4_1;
  wire bh40_w5_1;
  wire bh40_w6_1;
  wire bh40_w7_1;
  wire bh40_w8_1;
  wire bh40_w9_1;
  wire bh40_w10_1;
  wire bh40_w11_1;
  wire bh40_w12_1;
  wire bh40_w13_1;
  wire bh40_w14_1;
  wire bh40_w15_1;
  wire bh40_w16_1;
  wire bh40_w17_1;
  wire bh40_w18_1;
  wire bh40_w19_1;
  wire bh40_w20_1;
  wire bh40_w21_1;
  wire bh40_w22_1;
  wire bh40_w23_1;
  wire [28:0] bitheapfinaladd_bh40_in0;
  wire [28:0] bitheapfinaladd_bh40_in1;
  wire bitheapfinaladd_bh40_cin;
  wire [28:0] bitheapfinaladd_bh40_out;
  wire [28:0] bitheapresult_bh40;
  wire [28:0] outres;
  wire [4:0] n2216;
  wire [28:0] fixrealkcm_freq500_uid39_table0_n2217;
  wire n2220;
  wire n2221;
  wire n2222;
  wire n2223;
  wire n2224;
  wire n2225;
  wire n2226;
  wire n2227;
  wire n2228;
  wire n2229;
  wire n2230;
  wire n2231;
  wire n2232;
  wire n2233;
  wire n2234;
  wire n2235;
  wire n2236;
  wire n2237;
  wire n2238;
  wire n2239;
  wire n2240;
  wire n2241;
  wire n2242;
  wire n2243;
  wire n2244;
  wire n2245;
  wire n2246;
  wire n2247;
  wire n2248;
  wire [2:0] n2249;
  wire [23:0] fixrealkcm_freq500_uid39_table1_n2250;
  wire n2253;
  wire n2254;
  wire n2255;
  wire n2256;
  wire n2257;
  wire n2258;
  wire n2259;
  wire n2260;
  wire n2261;
  wire n2262;
  wire n2263;
  wire n2264;
  wire n2265;
  wire n2266;
  wire n2267;
  wire n2268;
  wire n2269;
  wire n2270;
  wire n2271;
  wire n2272;
  wire n2273;
  wire n2274;
  wire n2275;
  wire n2276;
  wire [1:0] n2278;
  wire [2:0] n2279;
  wire [3:0] n2280;
  wire [4:0] n2281;
  wire [5:0] n2282;
  wire [6:0] n2283;
  wire [7:0] n2284;
  wire [8:0] n2285;
  wire [9:0] n2286;
  wire [10:0] n2287;
  wire [11:0] n2288;
  wire [12:0] n2289;
  wire [13:0] n2290;
  wire [14:0] n2291;
  wire [15:0] n2292;
  wire [16:0] n2293;
  wire [17:0] n2294;
  wire [18:0] n2295;
  wire [19:0] n2296;
  wire [20:0] n2297;
  wire [21:0] n2298;
  wire [22:0] n2299;
  wire [23:0] n2300;
  wire [24:0] n2301;
  wire [25:0] n2302;
  wire [26:0] n2303;
  wire [27:0] n2304;
  wire [28:0] n2305;
  wire [5:0] n2307;
  wire [6:0] n2308;
  wire [7:0] n2309;
  wire [8:0] n2310;
  wire [9:0] n2311;
  wire [10:0] n2312;
  wire [11:0] n2313;
  wire [12:0] n2314;
  wire [13:0] n2315;
  wire [14:0] n2316;
  wire [15:0] n2317;
  wire [16:0] n2318;
  wire [17:0] n2319;
  wire [18:0] n2320;
  wire [19:0] n2321;
  wire [20:0] n2322;
  wire [21:0] n2323;
  wire [22:0] n2324;
  wire [23:0] n2325;
  wire [24:0] n2326;
  wire [25:0] n2327;
  wire [26:0] n2328;
  wire [27:0] n2329;
  wire [28:0] n2330;
  wire [28:0] bitheapfinaladd_bh40_n2332;
  reg [28:0] n2335;
  reg [23:0] n2336;
  assign r = outres; //(module output)
  /* fppowbf16.vhdl:2508:8  */
  assign fixrealkcm_freq500_uid39_a0 = n2216; // (signal)
  /* fppowbf16.vhdl:2510:8  */
  assign fixrealkcm_freq500_uid39_t0 = fixrealkcm_freq500_uid39_t0_copy43_d1; // (signal)
  /* fppowbf16.vhdl:2512:8  */
  assign fixrealkcm_freq500_uid39_t0_copy43 = fixrealkcm_freq500_uid39_table0_n2217; // (signal)
  /* fppowbf16.vhdl:2512:44  */
  assign fixrealkcm_freq500_uid39_t0_copy43_d1 = n2335; // (signal)
  /* fppowbf16.vhdl:2514:8  */
  assign bh40_w0_0 = n2220; // (signal)
  /* fppowbf16.vhdl:2516:8  */
  assign bh40_w1_0 = n2221; // (signal)
  /* fppowbf16.vhdl:2518:8  */
  assign bh40_w2_0 = n2222; // (signal)
  /* fppowbf16.vhdl:2520:8  */
  assign bh40_w3_0 = n2223; // (signal)
  /* fppowbf16.vhdl:2522:8  */
  assign bh40_w4_0 = n2224; // (signal)
  /* fppowbf16.vhdl:2524:8  */
  assign bh40_w5_0 = n2225; // (signal)
  /* fppowbf16.vhdl:2526:8  */
  assign bh40_w6_0 = n2226; // (signal)
  /* fppowbf16.vhdl:2528:8  */
  assign bh40_w7_0 = n2227; // (signal)
  /* fppowbf16.vhdl:2530:8  */
  assign bh40_w8_0 = n2228; // (signal)
  /* fppowbf16.vhdl:2532:8  */
  assign bh40_w9_0 = n2229; // (signal)
  /* fppowbf16.vhdl:2534:8  */
  assign bh40_w10_0 = n2230; // (signal)
  /* fppowbf16.vhdl:2536:8  */
  assign bh40_w11_0 = n2231; // (signal)
  /* fppowbf16.vhdl:2538:8  */
  assign bh40_w12_0 = n2232; // (signal)
  /* fppowbf16.vhdl:2540:8  */
  assign bh40_w13_0 = n2233; // (signal)
  /* fppowbf16.vhdl:2542:8  */
  assign bh40_w14_0 = n2234; // (signal)
  /* fppowbf16.vhdl:2544:8  */
  assign bh40_w15_0 = n2235; // (signal)
  /* fppowbf16.vhdl:2546:8  */
  assign bh40_w16_0 = n2236; // (signal)
  /* fppowbf16.vhdl:2548:8  */
  assign bh40_w17_0 = n2237; // (signal)
  /* fppowbf16.vhdl:2550:8  */
  assign bh40_w18_0 = n2238; // (signal)
  /* fppowbf16.vhdl:2552:8  */
  assign bh40_w19_0 = n2239; // (signal)
  /* fppowbf16.vhdl:2554:8  */
  assign bh40_w20_0 = n2240; // (signal)
  /* fppowbf16.vhdl:2556:8  */
  assign bh40_w21_0 = n2241; // (signal)
  /* fppowbf16.vhdl:2558:8  */
  assign bh40_w22_0 = n2242; // (signal)
  /* fppowbf16.vhdl:2560:8  */
  assign bh40_w23_0 = n2243; // (signal)
  /* fppowbf16.vhdl:2562:8  */
  assign bh40_w24_0 = n2244; // (signal)
  /* fppowbf16.vhdl:2564:8  */
  assign bh40_w25_0 = n2245; // (signal)
  /* fppowbf16.vhdl:2566:8  */
  assign bh40_w26_0 = n2246; // (signal)
  /* fppowbf16.vhdl:2568:8  */
  assign bh40_w27_0 = n2247; // (signal)
  /* fppowbf16.vhdl:2715:35  */
  assign bh40_w28_0 = n2248; // (signal)
  /* fppowbf16.vhdl:2572:8  */
  assign fixrealkcm_freq500_uid39_a1 = n2249; // (signal)
  /* fppowbf16.vhdl:2574:8  */
  assign fixrealkcm_freq500_uid39_t1 = fixrealkcm_freq500_uid39_t1_copy46_d1; // (signal)
  /* fppowbf16.vhdl:2576:8  */
  assign fixrealkcm_freq500_uid39_t1_copy46 = fixrealkcm_freq500_uid39_table1_n2250; // (signal)
  /* fppowbf16.vhdl:2576:44  */
  assign fixrealkcm_freq500_uid39_t1_copy46_d1 = n2336; // (signal)
  /* fppowbf16.vhdl:2578:8  */
  assign bh40_w0_1 = n2253; // (signal)
  /* fppowbf16.vhdl:2580:8  */
  assign bh40_w1_1 = n2254; // (signal)
  /* fppowbf16.vhdl:2582:8  */
  assign bh40_w2_1 = n2255; // (signal)
  /* fppowbf16.vhdl:2584:8  */
  assign bh40_w3_1 = n2256; // (signal)
  /* fppowbf16.vhdl:2586:8  */
  assign bh40_w4_1 = n2257; // (signal)
  /* fppowbf16.vhdl:2588:8  */
  assign bh40_w5_1 = n2258; // (signal)
  /* fppowbf16.vhdl:2590:8  */
  assign bh40_w6_1 = n2259; // (signal)
  /* fppowbf16.vhdl:2592:8  */
  assign bh40_w7_1 = n2260; // (signal)
  /* fppowbf16.vhdl:2594:8  */
  assign bh40_w8_1 = n2261; // (signal)
  /* fppowbf16.vhdl:2596:8  */
  assign bh40_w9_1 = n2262; // (signal)
  /* fppowbf16.vhdl:2598:8  */
  assign bh40_w10_1 = n2263; // (signal)
  /* fppowbf16.vhdl:2600:8  */
  assign bh40_w11_1 = n2264; // (signal)
  /* fppowbf16.vhdl:2602:8  */
  assign bh40_w12_1 = n2265; // (signal)
  /* fppowbf16.vhdl:2604:8  */
  assign bh40_w13_1 = n2266; // (signal)
  /* fppowbf16.vhdl:2606:8  */
  assign bh40_w14_1 = n2267; // (signal)
  /* fppowbf16.vhdl:2608:8  */
  assign bh40_w15_1 = n2268; // (signal)
  /* fppowbf16.vhdl:2610:8  */
  assign bh40_w16_1 = n2269; // (signal)
  /* fppowbf16.vhdl:2612:8  */
  assign bh40_w17_1 = n2270; // (signal)
  /* fppowbf16.vhdl:2614:8  */
  assign bh40_w18_1 = n2271; // (signal)
  /* fppowbf16.vhdl:2616:8  */
  assign bh40_w19_1 = n2272; // (signal)
  /* fppowbf16.vhdl:2618:8  */
  assign bh40_w20_1 = n2273; // (signal)
  /* fppowbf16.vhdl:2620:8  */
  assign bh40_w21_1 = n2274; // (signal)
  /* fppowbf16.vhdl:2622:8  */
  assign bh40_w22_1 = n2275; // (signal)
  /* fppowbf16.vhdl:2624:8  */
  assign bh40_w23_1 = n2276; // (signal)
  /* fppowbf16.vhdl:2626:8  */
  assign bitheapfinaladd_bh40_in0 = n2305; // (signal)
  /* fppowbf16.vhdl:2628:8  */
  assign bitheapfinaladd_bh40_in1 = n2330; // (signal)
  /* fppowbf16.vhdl:2630:8  */
  assign bitheapfinaladd_bh40_cin = 1'b0; // (signal)
  /* fppowbf16.vhdl:2632:8  */
  assign bitheapfinaladd_bh40_out = bitheapfinaladd_bh40_n2332; // (signal)
  /* fppowbf16.vhdl:2634:8  */
  assign bitheapresult_bh40 = bitheapfinaladd_bh40_out; // (signal)
  /* fppowbf16.vhdl:2636:8  */
  assign outres = bitheapresult_bh40; // (signal)
  /* fppowbf16.vhdl:2647:36  */
  assign n2216 = x[7:3]; // extract
  /* fppowbf16.vhdl:2648:4  */
  fixrealkcm_freq500_uid39_t0_freq500_uid42 fixrealkcm_freq500_uid39_table0 (
    .x(fixrealkcm_freq500_uid39_a0),
    .y(fixrealkcm_freq500_uid39_table0_n2217));
  /* fppowbf16.vhdl:2652:44  */
  assign n2220 = fixrealkcm_freq500_uid39_t0[0]; // extract
  /* fppowbf16.vhdl:2653:44  */
  assign n2221 = fixrealkcm_freq500_uid39_t0[1]; // extract
  /* fppowbf16.vhdl:2654:44  */
  assign n2222 = fixrealkcm_freq500_uid39_t0[2]; // extract
  /* fppowbf16.vhdl:2655:44  */
  assign n2223 = fixrealkcm_freq500_uid39_t0[3]; // extract
  /* fppowbf16.vhdl:2656:44  */
  assign n2224 = fixrealkcm_freq500_uid39_t0[4]; // extract
  /* fppowbf16.vhdl:2657:44  */
  assign n2225 = fixrealkcm_freq500_uid39_t0[5]; // extract
  /* fppowbf16.vhdl:2658:44  */
  assign n2226 = fixrealkcm_freq500_uid39_t0[6]; // extract
  /* fppowbf16.vhdl:2659:44  */
  assign n2227 = fixrealkcm_freq500_uid39_t0[7]; // extract
  /* fppowbf16.vhdl:2660:44  */
  assign n2228 = fixrealkcm_freq500_uid39_t0[8]; // extract
  /* fppowbf16.vhdl:2661:44  */
  assign n2229 = fixrealkcm_freq500_uid39_t0[9]; // extract
  /* fppowbf16.vhdl:2662:45  */
  assign n2230 = fixrealkcm_freq500_uid39_t0[10]; // extract
  /* fppowbf16.vhdl:2663:45  */
  assign n2231 = fixrealkcm_freq500_uid39_t0[11]; // extract
  /* fppowbf16.vhdl:2664:45  */
  assign n2232 = fixrealkcm_freq500_uid39_t0[12]; // extract
  /* fppowbf16.vhdl:2665:45  */
  assign n2233 = fixrealkcm_freq500_uid39_t0[13]; // extract
  /* fppowbf16.vhdl:2666:45  */
  assign n2234 = fixrealkcm_freq500_uid39_t0[14]; // extract
  /* fppowbf16.vhdl:2667:45  */
  assign n2235 = fixrealkcm_freq500_uid39_t0[15]; // extract
  /* fppowbf16.vhdl:2668:45  */
  assign n2236 = fixrealkcm_freq500_uid39_t0[16]; // extract
  /* fppowbf16.vhdl:2669:45  */
  assign n2237 = fixrealkcm_freq500_uid39_t0[17]; // extract
  /* fppowbf16.vhdl:2670:45  */
  assign n2238 = fixrealkcm_freq500_uid39_t0[18]; // extract
  /* fppowbf16.vhdl:2671:45  */
  assign n2239 = fixrealkcm_freq500_uid39_t0[19]; // extract
  /* fppowbf16.vhdl:2672:45  */
  assign n2240 = fixrealkcm_freq500_uid39_t0[20]; // extract
  /* fppowbf16.vhdl:2673:45  */
  assign n2241 = fixrealkcm_freq500_uid39_t0[21]; // extract
  /* fppowbf16.vhdl:2674:45  */
  assign n2242 = fixrealkcm_freq500_uid39_t0[22]; // extract
  /* fppowbf16.vhdl:2675:45  */
  assign n2243 = fixrealkcm_freq500_uid39_t0[23]; // extract
  /* fppowbf16.vhdl:2676:45  */
  assign n2244 = fixrealkcm_freq500_uid39_t0[24]; // extract
  /* fppowbf16.vhdl:2677:45  */
  assign n2245 = fixrealkcm_freq500_uid39_t0[25]; // extract
  /* fppowbf16.vhdl:2678:45  */
  assign n2246 = fixrealkcm_freq500_uid39_t0[26]; // extract
  /* fppowbf16.vhdl:2679:45  */
  assign n2247 = fixrealkcm_freq500_uid39_t0[27]; // extract
  /* fppowbf16.vhdl:2680:45  */
  assign n2248 = fixrealkcm_freq500_uid39_t0[28]; // extract
  /* fppowbf16.vhdl:2681:36  */
  assign n2249 = x[2:0]; // extract
  /* fppowbf16.vhdl:2682:4  */
  fixrealkcm_freq500_uid39_t1_freq500_uid45 fixrealkcm_freq500_uid39_table1 (
    .x(fixrealkcm_freq500_uid39_a1),
    .y(fixrealkcm_freq500_uid39_table1_n2250));
  /* fppowbf16.vhdl:2686:44  */
  assign n2253 = fixrealkcm_freq500_uid39_t1[0]; // extract
  /* fppowbf16.vhdl:2687:44  */
  assign n2254 = fixrealkcm_freq500_uid39_t1[1]; // extract
  /* fppowbf16.vhdl:2688:44  */
  assign n2255 = fixrealkcm_freq500_uid39_t1[2]; // extract
  /* fppowbf16.vhdl:2689:44  */
  assign n2256 = fixrealkcm_freq500_uid39_t1[3]; // extract
  /* fppowbf16.vhdl:2690:44  */
  assign n2257 = fixrealkcm_freq500_uid39_t1[4]; // extract
  /* fppowbf16.vhdl:2691:44  */
  assign n2258 = fixrealkcm_freq500_uid39_t1[5]; // extract
  /* fppowbf16.vhdl:2692:44  */
  assign n2259 = fixrealkcm_freq500_uid39_t1[6]; // extract
  /* fppowbf16.vhdl:2693:44  */
  assign n2260 = fixrealkcm_freq500_uid39_t1[7]; // extract
  /* fppowbf16.vhdl:2694:44  */
  assign n2261 = fixrealkcm_freq500_uid39_t1[8]; // extract
  /* fppowbf16.vhdl:2695:44  */
  assign n2262 = fixrealkcm_freq500_uid39_t1[9]; // extract
  /* fppowbf16.vhdl:2696:45  */
  assign n2263 = fixrealkcm_freq500_uid39_t1[10]; // extract
  /* fppowbf16.vhdl:2697:45  */
  assign n2264 = fixrealkcm_freq500_uid39_t1[11]; // extract
  /* fppowbf16.vhdl:2698:45  */
  assign n2265 = fixrealkcm_freq500_uid39_t1[12]; // extract
  /* fppowbf16.vhdl:2699:45  */
  assign n2266 = fixrealkcm_freq500_uid39_t1[13]; // extract
  /* fppowbf16.vhdl:2700:45  */
  assign n2267 = fixrealkcm_freq500_uid39_t1[14]; // extract
  /* fppowbf16.vhdl:2701:45  */
  assign n2268 = fixrealkcm_freq500_uid39_t1[15]; // extract
  /* fppowbf16.vhdl:2702:45  */
  assign n2269 = fixrealkcm_freq500_uid39_t1[16]; // extract
  /* fppowbf16.vhdl:2703:45  */
  assign n2270 = fixrealkcm_freq500_uid39_t1[17]; // extract
  /* fppowbf16.vhdl:2704:45  */
  assign n2271 = fixrealkcm_freq500_uid39_t1[18]; // extract
  /* fppowbf16.vhdl:2705:45  */
  assign n2272 = fixrealkcm_freq500_uid39_t1[19]; // extract
  /* fppowbf16.vhdl:2706:45  */
  assign n2273 = fixrealkcm_freq500_uid39_t1[20]; // extract
  /* fppowbf16.vhdl:2707:45  */
  assign n2274 = fixrealkcm_freq500_uid39_t1[21]; // extract
  /* fppowbf16.vhdl:2708:45  */
  assign n2275 = fixrealkcm_freq500_uid39_t1[22]; // extract
  /* fppowbf16.vhdl:2709:45  */
  assign n2276 = fixrealkcm_freq500_uid39_t1[23]; // extract
  /* fppowbf16.vhdl:2715:48  */
  assign n2278 = {bh40_w28_0, bh40_w27_0};
  /* fppowbf16.vhdl:2715:61  */
  assign n2279 = {n2278, bh40_w26_0};
  /* fppowbf16.vhdl:2715:74  */
  assign n2280 = {n2279, bh40_w25_0};
  /* fppowbf16.vhdl:2715:87  */
  assign n2281 = {n2280, bh40_w24_0};
  /* fppowbf16.vhdl:2715:100  */
  assign n2282 = {n2281, bh40_w23_1};
  /* fppowbf16.vhdl:2715:113  */
  assign n2283 = {n2282, bh40_w22_1};
  /* fppowbf16.vhdl:2715:126  */
  assign n2284 = {n2283, bh40_w21_1};
  /* fppowbf16.vhdl:2715:139  */
  assign n2285 = {n2284, bh40_w20_1};
  /* fppowbf16.vhdl:2715:152  */
  assign n2286 = {n2285, bh40_w19_1};
  /* fppowbf16.vhdl:2715:165  */
  assign n2287 = {n2286, bh40_w18_1};
  /* fppowbf16.vhdl:2715:178  */
  assign n2288 = {n2287, bh40_w17_1};
  /* fppowbf16.vhdl:2715:191  */
  assign n2289 = {n2288, bh40_w16_1};
  /* fppowbf16.vhdl:2715:204  */
  assign n2290 = {n2289, bh40_w15_1};
  /* fppowbf16.vhdl:2715:217  */
  assign n2291 = {n2290, bh40_w14_1};
  /* fppowbf16.vhdl:2715:230  */
  assign n2292 = {n2291, bh40_w13_1};
  /* fppowbf16.vhdl:2715:243  */
  assign n2293 = {n2292, bh40_w12_1};
  /* fppowbf16.vhdl:2715:256  */
  assign n2294 = {n2293, bh40_w11_1};
  /* fppowbf16.vhdl:2715:269  */
  assign n2295 = {n2294, bh40_w10_1};
  /* fppowbf16.vhdl:2715:282  */
  assign n2296 = {n2295, bh40_w9_1};
  /* fppowbf16.vhdl:2715:294  */
  assign n2297 = {n2296, bh40_w8_1};
  /* fppowbf16.vhdl:2715:306  */
  assign n2298 = {n2297, bh40_w7_1};
  /* fppowbf16.vhdl:2715:318  */
  assign n2299 = {n2298, bh40_w6_1};
  /* fppowbf16.vhdl:2715:330  */
  assign n2300 = {n2299, bh40_w5_1};
  /* fppowbf16.vhdl:2715:342  */
  assign n2301 = {n2300, bh40_w4_1};
  /* fppowbf16.vhdl:2715:354  */
  assign n2302 = {n2301, bh40_w3_1};
  /* fppowbf16.vhdl:2715:366  */
  assign n2303 = {n2302, bh40_w2_1};
  /* fppowbf16.vhdl:2715:378  */
  assign n2304 = {n2303, bh40_w1_1};
  /* fppowbf16.vhdl:2715:390  */
  assign n2305 = {n2304, bh40_w0_1};
  /* fppowbf16.vhdl:2716:60  */
  assign n2307 = {5'b00000, bh40_w23_0};
  /* fppowbf16.vhdl:2716:73  */
  assign n2308 = {n2307, bh40_w22_0};
  /* fppowbf16.vhdl:2716:86  */
  assign n2309 = {n2308, bh40_w21_0};
  /* fppowbf16.vhdl:2716:99  */
  assign n2310 = {n2309, bh40_w20_0};
  /* fppowbf16.vhdl:2716:112  */
  assign n2311 = {n2310, bh40_w19_0};
  /* fppowbf16.vhdl:2716:125  */
  assign n2312 = {n2311, bh40_w18_0};
  /* fppowbf16.vhdl:2716:138  */
  assign n2313 = {n2312, bh40_w17_0};
  /* fppowbf16.vhdl:2716:151  */
  assign n2314 = {n2313, bh40_w16_0};
  /* fppowbf16.vhdl:2716:164  */
  assign n2315 = {n2314, bh40_w15_0};
  /* fppowbf16.vhdl:2716:177  */
  assign n2316 = {n2315, bh40_w14_0};
  /* fppowbf16.vhdl:2716:190  */
  assign n2317 = {n2316, bh40_w13_0};
  /* fppowbf16.vhdl:2716:203  */
  assign n2318 = {n2317, bh40_w12_0};
  /* fppowbf16.vhdl:2716:216  */
  assign n2319 = {n2318, bh40_w11_0};
  /* fppowbf16.vhdl:2716:229  */
  assign n2320 = {n2319, bh40_w10_0};
  /* fppowbf16.vhdl:2716:242  */
  assign n2321 = {n2320, bh40_w9_0};
  /* fppowbf16.vhdl:2716:254  */
  assign n2322 = {n2321, bh40_w8_0};
  /* fppowbf16.vhdl:2716:266  */
  assign n2323 = {n2322, bh40_w7_0};
  /* fppowbf16.vhdl:2716:278  */
  assign n2324 = {n2323, bh40_w6_0};
  /* fppowbf16.vhdl:2716:290  */
  assign n2325 = {n2324, bh40_w5_0};
  /* fppowbf16.vhdl:2716:302  */
  assign n2326 = {n2325, bh40_w4_0};
  /* fppowbf16.vhdl:2716:314  */
  assign n2327 = {n2326, bh40_w3_0};
  /* fppowbf16.vhdl:2716:326  */
  assign n2328 = {n2327, bh40_w2_0};
  /* fppowbf16.vhdl:2716:338  */
  assign n2329 = {n2328, bh40_w1_0};
  /* fppowbf16.vhdl:2716:350  */
  assign n2330 = {n2329, bh40_w0_0};
  /* fppowbf16.vhdl:2719:4  */
  intadder_29_freq500_uid49 bitheapfinaladd_bh40 (
    .clk(clk),
    .x(bitheapfinaladd_bh40_in0),
    .y(bitheapfinaladd_bh40_in1),
    .cin(bitheapfinaladd_bh40_cin),
    .r(bitheapfinaladd_bh40_n2332));
  /* fppowbf16.vhdl:2641:10  */
  always @(posedge clk)
    n2335 <= fixrealkcm_freq500_uid39_t0_copy43;
  /* fppowbf16.vhdl:2641:10  */
  always @(posedge clk)
    n2336 <= fixrealkcm_freq500_uid39_t1_copy46;
endmodule

module intadder_30_freq500_uid37
  (input  clk,
   input  [29:0] x,
   input  [29:0] y,
   input  cin,
   output [29:0] r);
  wire [29:0] rtmp;
  wire [29:0] x_d1;
  wire [29:0] x_d2;
  wire [29:0] x_d3;
  wire [29:0] x_d4;
  wire cin_d1;
  wire cin_d2;
  wire cin_d3;
  wire cin_d4;
  wire cin_d5;
  wire cin_d6;
  wire [29:0] n2196;
  wire [29:0] n2197;
  wire [29:0] n2198;
  reg [29:0] n2199;
  reg [29:0] n2200;
  reg [29:0] n2201;
  reg [29:0] n2202;
  reg n2203;
  reg n2204;
  reg n2205;
  reg n2206;
  reg n2207;
  reg n2208;
  assign r = rtmp; //(module output)
  /* fppowbf16.vhdl:2387:8  */
  assign rtmp = n2198; // (signal)
  /* fppowbf16.vhdl:2389:8  */
  assign x_d1 = n2199; // (signal)
  /* fppowbf16.vhdl:2389:14  */
  assign x_d2 = n2200; // (signal)
  /* fppowbf16.vhdl:2389:20  */
  assign x_d3 = n2201; // (signal)
  /* fppowbf16.vhdl:2389:26  */
  assign x_d4 = n2202; // (signal)
  /* fppowbf16.vhdl:2391:8  */
  assign cin_d1 = n2203; // (signal)
  /* fppowbf16.vhdl:2391:16  */
  assign cin_d2 = n2204; // (signal)
  /* fppowbf16.vhdl:2391:24  */
  assign cin_d3 = n2205; // (signal)
  /* fppowbf16.vhdl:2391:32  */
  assign cin_d4 = n2206; // (signal)
  /* fppowbf16.vhdl:2391:40  */
  assign cin_d5 = n2207; // (signal)
  /* fppowbf16.vhdl:2391:48  */
  assign cin_d6 = n2208; // (signal)
  /* fppowbf16.vhdl:2409:17  */
  assign n2196 = x_d4 + y;
  /* fppowbf16.vhdl:2409:21  */
  assign n2197 = {29'b0, cin_d6};  //  uext
  /* fppowbf16.vhdl:2409:21  */
  assign n2198 = n2196 + n2197;
  /* fppowbf16.vhdl:2396:10  */
  always @(posedge clk)
    n2199 <= x;
  /* fppowbf16.vhdl:2396:10  */
  always @(posedge clk)
    n2200 <= x_d1;
  /* fppowbf16.vhdl:2396:10  */
  always @(posedge clk)
    n2201 <= x_d2;
  /* fppowbf16.vhdl:2396:10  */
  always @(posedge clk)
    n2202 <= x_d3;
  /* fppowbf16.vhdl:2396:10  */
  always @(posedge clk)
    n2203 <= cin;
  /* fppowbf16.vhdl:2396:10  */
  always @(posedge clk)
    n2204 <= cin_d1;
  /* fppowbf16.vhdl:2396:10  */
  always @(posedge clk)
    n2205 <= cin_d2;
  /* fppowbf16.vhdl:2396:10  */
  always @(posedge clk)
    n2206 <= cin_d3;
  /* fppowbf16.vhdl:2396:10  */
  always @(posedge clk)
    n2207 <= cin_d4;
  /* fppowbf16.vhdl:2396:10  */
  always @(posedge clk)
    n2208 <= cin_d5;
endmodule

module intadder_30_freq500_uid34
  (input  clk,
   input  [29:0] x,
   input  [29:0] y,
   input  cin,
   output [29:0] r);
  wire cin_1;
  wire cin_1_d1;
  wire cin_1_d2;
  wire [30:0] x_1;
  wire [30:0] x_1_d1;
  wire [30:0] x_1_d2;
  wire [30:0] y_1;
  wire [30:0] y_1_d1;
  wire [30:0] s_1;
  wire [29:0] r_1;
  wire [30:0] n2169;
  wire [30:0] n2171;
  wire [30:0] n2172;
  wire [30:0] n2173;
  wire [30:0] n2174;
  wire [29:0] n2175;
  reg n2176;
  reg n2177;
  reg [30:0] n2178;
  reg [30:0] n2179;
  reg [30:0] n2180;
  assign r = r_1; //(module output)
  /* fppowbf16.vhdl:2326:15  */
  assign cin_1_d1 = n2176; // (signal)
  /* fppowbf16.vhdl:2326:25  */
  assign cin_1_d2 = n2177; // (signal)
  /* fppowbf16.vhdl:2328:8  */
  assign x_1 = n2169; // (signal)
  /* fppowbf16.vhdl:2328:13  */
  assign x_1_d1 = n2178; // (signal)
  /* fppowbf16.vhdl:2328:21  */
  assign x_1_d2 = n2179; // (signal)
  /* fppowbf16.vhdl:2330:8  */
  assign y_1 = n2171; // (signal)
  /* fppowbf16.vhdl:2330:13  */
  assign y_1_d1 = n2180; // (signal)
  /* fppowbf16.vhdl:2332:8  */
  assign s_1 = n2174; // (signal)
  /* fppowbf16.vhdl:2334:8  */
  assign r_1 = n2175; // (signal)
  /* fppowbf16.vhdl:2348:15  */
  assign n2169 = {1'b0, x};
  /* fppowbf16.vhdl:2349:15  */
  assign n2171 = {1'b0, y};
  /* fppowbf16.vhdl:2350:18  */
  assign n2172 = x_1_d2 + y_1_d1;
  /* fppowbf16.vhdl:2350:27  */
  assign n2173 = {30'b0, cin_1_d2};  //  uext
  /* fppowbf16.vhdl:2350:27  */
  assign n2174 = n2172 + n2173;
  /* fppowbf16.vhdl:2351:14  */
  assign n2175 = s_1[29:0]; // extract
  /* fppowbf16.vhdl:2339:10  */
  always @(posedge clk)
    n2176 <= cin_1;
  /* fppowbf16.vhdl:2339:10  */
  always @(posedge clk)
    n2177 <= cin_1_d1;
  /* fppowbf16.vhdl:2339:10  */
  always @(posedge clk)
    n2178 <= x_1;
  /* fppowbf16.vhdl:2339:10  */
  always @(posedge clk)
    n2179 <= x_1_d1;
  /* fppowbf16.vhdl:2339:10  */
  always @(posedge clk)
    n2180 <= y_1;
endmodule

module logtable1_freq500_uid30
  (input  [4:0] x,
   output [24:0] y);
  wire [24:0] y0;
  wire [24:0] y1;
  wire n2061;
  wire n2064;
  wire n2067;
  wire n2070;
  wire n2073;
  wire n2076;
  wire n2079;
  wire n2082;
  wire n2085;
  wire n2088;
  wire n2091;
  wire n2094;
  wire n2097;
  wire n2100;
  wire n2103;
  wire n2106;
  wire n2109;
  wire n2112;
  wire n2115;
  wire n2118;
  wire n2121;
  wire n2124;
  wire n2127;
  wire n2130;
  wire n2133;
  wire n2136;
  wire n2139;
  wire n2142;
  wire n2145;
  wire n2148;
  wire n2151;
  wire n2154;
  wire [31:0] n2156;
  reg [24:0] n2157;
  assign y = y1; //(module output)
  /* fppowbf16.vhdl:366:8  */
  assign y0 = n2157; // (signal)
  /* fppowbf16.vhdl:368:8  */
  assign y1 = y0; // (signal)
  /* fppowbf16.vhdl:372:35  */
  assign n2061 = x == 5'b00000;
  /* fppowbf16.vhdl:373:35  */
  assign n2064 = x == 5'b00001;
  /* fppowbf16.vhdl:374:35  */
  assign n2067 = x == 5'b00010;
  /* fppowbf16.vhdl:375:35  */
  assign n2070 = x == 5'b00011;
  /* fppowbf16.vhdl:376:35  */
  assign n2073 = x == 5'b00100;
  /* fppowbf16.vhdl:377:35  */
  assign n2076 = x == 5'b00101;
  /* fppowbf16.vhdl:378:35  */
  assign n2079 = x == 5'b00110;
  /* fppowbf16.vhdl:379:35  */
  assign n2082 = x == 5'b00111;
  /* fppowbf16.vhdl:380:35  */
  assign n2085 = x == 5'b01000;
  /* fppowbf16.vhdl:381:35  */
  assign n2088 = x == 5'b01001;
  /* fppowbf16.vhdl:382:35  */
  assign n2091 = x == 5'b01010;
  /* fppowbf16.vhdl:383:35  */
  assign n2094 = x == 5'b01011;
  /* fppowbf16.vhdl:384:35  */
  assign n2097 = x == 5'b01100;
  /* fppowbf16.vhdl:385:35  */
  assign n2100 = x == 5'b01101;
  /* fppowbf16.vhdl:386:35  */
  assign n2103 = x == 5'b01110;
  /* fppowbf16.vhdl:387:35  */
  assign n2106 = x == 5'b01111;
  /* fppowbf16.vhdl:388:35  */
  assign n2109 = x == 5'b10000;
  /* fppowbf16.vhdl:389:35  */
  assign n2112 = x == 5'b10001;
  /* fppowbf16.vhdl:390:35  */
  assign n2115 = x == 5'b10010;
  /* fppowbf16.vhdl:391:35  */
  assign n2118 = x == 5'b10011;
  /* fppowbf16.vhdl:392:35  */
  assign n2121 = x == 5'b10100;
  /* fppowbf16.vhdl:393:35  */
  assign n2124 = x == 5'b10101;
  /* fppowbf16.vhdl:394:35  */
  assign n2127 = x == 5'b10110;
  /* fppowbf16.vhdl:395:35  */
  assign n2130 = x == 5'b10111;
  /* fppowbf16.vhdl:396:35  */
  assign n2133 = x == 5'b11000;
  /* fppowbf16.vhdl:397:35  */
  assign n2136 = x == 5'b11001;
  /* fppowbf16.vhdl:398:35  */
  assign n2139 = x == 5'b11010;
  /* fppowbf16.vhdl:399:35  */
  assign n2142 = x == 5'b11011;
  /* fppowbf16.vhdl:400:35  */
  assign n2145 = x == 5'b11100;
  /* fppowbf16.vhdl:401:35  */
  assign n2148 = x == 5'b11101;
  /* fppowbf16.vhdl:402:35  */
  assign n2151 = x == 5'b11110;
  /* fppowbf16.vhdl:403:35  */
  assign n2154 = x == 5'b11111;
  assign n2156 = {n2154, n2151, n2148, n2145, n2142, n2139, n2136, n2133, n2130, n2127, n2124, n2121, n2118, n2115, n2112, n2109, n2106, n2103, n2100, n2097, n2094, n2091, n2088, n2085, n2082, n2079, n2076, n2073, n2070, n2067, n2064, n2061};
  /* fppowbf16.vhdl:371:4  */
  always @*
    case (n2156)
      32'b10000000000000000000000000000000: n2157 = 25'b1111101110010101111110011;
      32'b01000000000000000000000000000000: n2157 = 25'b1111001101011001001110010;
      32'b00100000000000000000000000000000: n2157 = 25'b1110101100011110100101111;
      32'b00010000000000000000000000000000: n2157 = 25'b1110001011100110000100110;
      32'b00001000000000000000000000000000: n2157 = 25'b1101101010101111101010101;
      32'b00000100000000000000000000000000: n2157 = 25'b1101001001111011010111010;
      32'b00000010000000000000000000000000: n2157 = 25'b1100101001001001001010011;
      32'b00000001000000000000000000000000: n2157 = 25'b1100001000011001000011101;
      32'b00000000100000000000000000000000: n2157 = 25'b1011100111101011000011000;
      32'b00000000010000000000000000000000: n2157 = 25'b1011000110111111000111111;
      32'b00000000001000000000000000000000: n2157 = 25'b1010100110010101010010010;
      32'b00000000000100000000000000000000: n2157 = 25'b1010000101101101100001111;
      32'b00000000000010000000000000000000: n2157 = 25'b1001100101000111110110010;
      32'b00000000000001000000000000000000: n2157 = 25'b1001000100100100001111010;
      32'b00000000000000100000000000000000: n2157 = 25'b1000100100000010101100110;
      32'b00000000000000010000000000000000: n2157 = 25'b1000000011100011001110010;
      32'b00000000000000001000000000000000: n2157 = 25'b0111110011010100010000011;
      32'b00000000000000000100000000000000: n2157 = 25'b0111010010110111110111100;
      32'b00000000000000000010000000000000: n2157 = 25'b0110110010011101100010001;
      32'b00000000000000000001000000000000: n2157 = 25'b0110010010000101010000000;
      32'b00000000000000000000100000000000: n2157 = 25'b0101110001101111000000101;
      32'b00000000000000000000010000000000: n2157 = 25'b0101010001011010110100000;
      32'b00000000000000000000001000000000: n2157 = 25'b0100110001001000101001110;
      32'b00000000000000000000000100000000: n2157 = 25'b0100010000111000100001110;
      32'b00000000000000000000000010000000: n2157 = 25'b0011110000101010011011100;
      32'b00000000000000000000000001000000: n2157 = 25'b0011010000011110010111000;
      32'b00000000000000000000000000100000: n2157 = 25'b0010110000010100010011110;
      32'b00000000000000000000000000010000: n2157 = 25'b0010010000001100010001110;
      32'b00000000000000000000000000001000: n2157 = 25'b0001110000000110010000101;
      32'b00000000000000000000000000000100: n2157 = 25'b0001010000000010010000001;
      32'b00000000000000000000000000000010: n2157 = 25'b0000110000000000010000000;
      32'b00000000000000000000000000000001: n2157 = 25'b0000010000000000010000000;
      default: n2157 = 25'bX;
    endcase
endmodule

module logtable0_freq500_uid27
  (input  [6:0] x,
   output [29:0] y);
  wire [29:0] y0;
  wire [29:0] y1;
  wire n1673;
  wire n1676;
  wire n1679;
  wire n1682;
  wire n1685;
  wire n1688;
  wire n1691;
  wire n1694;
  wire n1697;
  wire n1700;
  wire n1703;
  wire n1706;
  wire n1709;
  wire n1712;
  wire n1715;
  wire n1718;
  wire n1721;
  wire n1724;
  wire n1727;
  wire n1730;
  wire n1733;
  wire n1736;
  wire n1739;
  wire n1742;
  wire n1745;
  wire n1748;
  wire n1751;
  wire n1754;
  wire n1757;
  wire n1760;
  wire n1763;
  wire n1766;
  wire n1769;
  wire n1772;
  wire n1775;
  wire n1778;
  wire n1781;
  wire n1784;
  wire n1787;
  wire n1790;
  wire n1793;
  wire n1796;
  wire n1799;
  wire n1802;
  wire n1805;
  wire n1808;
  wire n1811;
  wire n1814;
  wire n1817;
  wire n1820;
  wire n1823;
  wire n1826;
  wire n1829;
  wire n1832;
  wire n1835;
  wire n1838;
  wire n1841;
  wire n1844;
  wire n1847;
  wire n1850;
  wire n1853;
  wire n1856;
  wire n1859;
  wire n1862;
  wire n1865;
  wire n1868;
  wire n1871;
  wire n1874;
  wire n1877;
  wire n1880;
  wire n1883;
  wire n1886;
  wire n1889;
  wire n1892;
  wire n1895;
  wire n1898;
  wire n1901;
  wire n1904;
  wire n1907;
  wire n1910;
  wire n1913;
  wire n1916;
  wire n1919;
  wire n1922;
  wire n1925;
  wire n1928;
  wire n1931;
  wire n1934;
  wire n1937;
  wire n1940;
  wire n1943;
  wire n1946;
  wire n1949;
  wire n1952;
  wire n1955;
  wire n1958;
  wire n1961;
  wire n1964;
  wire n1967;
  wire n1970;
  wire n1973;
  wire n1976;
  wire n1979;
  wire n1982;
  wire n1985;
  wire n1988;
  wire n1991;
  wire n1994;
  wire n1997;
  wire n2000;
  wire n2003;
  wire n2006;
  wire n2009;
  wire n2012;
  wire n2015;
  wire n2018;
  wire n2021;
  wire n2024;
  wire n2027;
  wire n2030;
  wire n2033;
  wire n2036;
  wire n2039;
  wire n2042;
  wire n2045;
  wire n2048;
  wire n2051;
  wire n2054;
  wire [127:0] n2056;
  reg [29:0] n2057;
  assign y = y1; //(module output)
  /* fppowbf16.vhdl:198:8  */
  assign y0 = n2057; // (signal)
  /* fppowbf16.vhdl:200:8  */
  assign y1 = y0; // (signal)
  /* fppowbf16.vhdl:204:40  */
  assign n1673 = x == 7'b0000000;
  /* fppowbf16.vhdl:205:40  */
  assign n1676 = x == 7'b0000001;
  /* fppowbf16.vhdl:206:40  */
  assign n1679 = x == 7'b0000010;
  /* fppowbf16.vhdl:207:40  */
  assign n1682 = x == 7'b0000011;
  /* fppowbf16.vhdl:208:40  */
  assign n1685 = x == 7'b0000100;
  /* fppowbf16.vhdl:209:40  */
  assign n1688 = x == 7'b0000101;
  /* fppowbf16.vhdl:210:40  */
  assign n1691 = x == 7'b0000110;
  /* fppowbf16.vhdl:211:40  */
  assign n1694 = x == 7'b0000111;
  /* fppowbf16.vhdl:212:40  */
  assign n1697 = x == 7'b0001000;
  /* fppowbf16.vhdl:213:40  */
  assign n1700 = x == 7'b0001001;
  /* fppowbf16.vhdl:214:40  */
  assign n1703 = x == 7'b0001010;
  /* fppowbf16.vhdl:215:40  */
  assign n1706 = x == 7'b0001011;
  /* fppowbf16.vhdl:216:40  */
  assign n1709 = x == 7'b0001100;
  /* fppowbf16.vhdl:217:40  */
  assign n1712 = x == 7'b0001101;
  /* fppowbf16.vhdl:218:40  */
  assign n1715 = x == 7'b0001110;
  /* fppowbf16.vhdl:219:40  */
  assign n1718 = x == 7'b0001111;
  /* fppowbf16.vhdl:220:40  */
  assign n1721 = x == 7'b0010000;
  /* fppowbf16.vhdl:221:40  */
  assign n1724 = x == 7'b0010001;
  /* fppowbf16.vhdl:222:40  */
  assign n1727 = x == 7'b0010010;
  /* fppowbf16.vhdl:223:40  */
  assign n1730 = x == 7'b0010011;
  /* fppowbf16.vhdl:224:40  */
  assign n1733 = x == 7'b0010100;
  /* fppowbf16.vhdl:225:40  */
  assign n1736 = x == 7'b0010101;
  /* fppowbf16.vhdl:226:40  */
  assign n1739 = x == 7'b0010110;
  /* fppowbf16.vhdl:227:40  */
  assign n1742 = x == 7'b0010111;
  /* fppowbf16.vhdl:228:40  */
  assign n1745 = x == 7'b0011000;
  /* fppowbf16.vhdl:229:40  */
  assign n1748 = x == 7'b0011001;
  /* fppowbf16.vhdl:230:40  */
  assign n1751 = x == 7'b0011010;
  /* fppowbf16.vhdl:231:40  */
  assign n1754 = x == 7'b0011011;
  /* fppowbf16.vhdl:232:40  */
  assign n1757 = x == 7'b0011100;
  /* fppowbf16.vhdl:233:40  */
  assign n1760 = x == 7'b0011101;
  /* fppowbf16.vhdl:234:40  */
  assign n1763 = x == 7'b0011110;
  /* fppowbf16.vhdl:235:40  */
  assign n1766 = x == 7'b0011111;
  /* fppowbf16.vhdl:236:40  */
  assign n1769 = x == 7'b0100000;
  /* fppowbf16.vhdl:237:40  */
  assign n1772 = x == 7'b0100001;
  /* fppowbf16.vhdl:238:40  */
  assign n1775 = x == 7'b0100010;
  /* fppowbf16.vhdl:239:40  */
  assign n1778 = x == 7'b0100011;
  /* fppowbf16.vhdl:240:40  */
  assign n1781 = x == 7'b0100100;
  /* fppowbf16.vhdl:241:40  */
  assign n1784 = x == 7'b0100101;
  /* fppowbf16.vhdl:242:40  */
  assign n1787 = x == 7'b0100110;
  /* fppowbf16.vhdl:243:40  */
  assign n1790 = x == 7'b0100111;
  /* fppowbf16.vhdl:244:40  */
  assign n1793 = x == 7'b0101000;
  /* fppowbf16.vhdl:245:40  */
  assign n1796 = x == 7'b0101001;
  /* fppowbf16.vhdl:246:40  */
  assign n1799 = x == 7'b0101010;
  /* fppowbf16.vhdl:247:40  */
  assign n1802 = x == 7'b0101011;
  /* fppowbf16.vhdl:248:40  */
  assign n1805 = x == 7'b0101100;
  /* fppowbf16.vhdl:249:40  */
  assign n1808 = x == 7'b0101101;
  /* fppowbf16.vhdl:250:40  */
  assign n1811 = x == 7'b0101110;
  /* fppowbf16.vhdl:251:40  */
  assign n1814 = x == 7'b0101111;
  /* fppowbf16.vhdl:252:40  */
  assign n1817 = x == 7'b0110000;
  /* fppowbf16.vhdl:253:40  */
  assign n1820 = x == 7'b0110001;
  /* fppowbf16.vhdl:254:40  */
  assign n1823 = x == 7'b0110010;
  /* fppowbf16.vhdl:255:40  */
  assign n1826 = x == 7'b0110011;
  /* fppowbf16.vhdl:256:40  */
  assign n1829 = x == 7'b0110100;
  /* fppowbf16.vhdl:257:40  */
  assign n1832 = x == 7'b0110101;
  /* fppowbf16.vhdl:258:40  */
  assign n1835 = x == 7'b0110110;
  /* fppowbf16.vhdl:259:40  */
  assign n1838 = x == 7'b0110111;
  /* fppowbf16.vhdl:260:40  */
  assign n1841 = x == 7'b0111000;
  /* fppowbf16.vhdl:261:40  */
  assign n1844 = x == 7'b0111001;
  /* fppowbf16.vhdl:262:40  */
  assign n1847 = x == 7'b0111010;
  /* fppowbf16.vhdl:263:40  */
  assign n1850 = x == 7'b0111011;
  /* fppowbf16.vhdl:264:40  */
  assign n1853 = x == 7'b0111100;
  /* fppowbf16.vhdl:265:40  */
  assign n1856 = x == 7'b0111101;
  /* fppowbf16.vhdl:266:40  */
  assign n1859 = x == 7'b0111110;
  /* fppowbf16.vhdl:267:40  */
  assign n1862 = x == 7'b0111111;
  /* fppowbf16.vhdl:268:40  */
  assign n1865 = x == 7'b1000000;
  /* fppowbf16.vhdl:269:40  */
  assign n1868 = x == 7'b1000001;
  /* fppowbf16.vhdl:270:40  */
  assign n1871 = x == 7'b1000010;
  /* fppowbf16.vhdl:271:40  */
  assign n1874 = x == 7'b1000011;
  /* fppowbf16.vhdl:272:40  */
  assign n1877 = x == 7'b1000100;
  /* fppowbf16.vhdl:273:40  */
  assign n1880 = x == 7'b1000101;
  /* fppowbf16.vhdl:274:40  */
  assign n1883 = x == 7'b1000110;
  /* fppowbf16.vhdl:275:40  */
  assign n1886 = x == 7'b1000111;
  /* fppowbf16.vhdl:276:40  */
  assign n1889 = x == 7'b1001000;
  /* fppowbf16.vhdl:277:40  */
  assign n1892 = x == 7'b1001001;
  /* fppowbf16.vhdl:278:40  */
  assign n1895 = x == 7'b1001010;
  /* fppowbf16.vhdl:279:40  */
  assign n1898 = x == 7'b1001011;
  /* fppowbf16.vhdl:280:40  */
  assign n1901 = x == 7'b1001100;
  /* fppowbf16.vhdl:281:40  */
  assign n1904 = x == 7'b1001101;
  /* fppowbf16.vhdl:282:40  */
  assign n1907 = x == 7'b1001110;
  /* fppowbf16.vhdl:283:40  */
  assign n1910 = x == 7'b1001111;
  /* fppowbf16.vhdl:284:40  */
  assign n1913 = x == 7'b1010000;
  /* fppowbf16.vhdl:285:40  */
  assign n1916 = x == 7'b1010001;
  /* fppowbf16.vhdl:286:40  */
  assign n1919 = x == 7'b1010010;
  /* fppowbf16.vhdl:287:40  */
  assign n1922 = x == 7'b1010011;
  /* fppowbf16.vhdl:288:40  */
  assign n1925 = x == 7'b1010100;
  /* fppowbf16.vhdl:289:40  */
  assign n1928 = x == 7'b1010101;
  /* fppowbf16.vhdl:290:40  */
  assign n1931 = x == 7'b1010110;
  /* fppowbf16.vhdl:291:40  */
  assign n1934 = x == 7'b1010111;
  /* fppowbf16.vhdl:292:40  */
  assign n1937 = x == 7'b1011000;
  /* fppowbf16.vhdl:293:40  */
  assign n1940 = x == 7'b1011001;
  /* fppowbf16.vhdl:294:40  */
  assign n1943 = x == 7'b1011010;
  /* fppowbf16.vhdl:295:40  */
  assign n1946 = x == 7'b1011011;
  /* fppowbf16.vhdl:296:40  */
  assign n1949 = x == 7'b1011100;
  /* fppowbf16.vhdl:297:40  */
  assign n1952 = x == 7'b1011101;
  /* fppowbf16.vhdl:298:40  */
  assign n1955 = x == 7'b1011110;
  /* fppowbf16.vhdl:299:40  */
  assign n1958 = x == 7'b1011111;
  /* fppowbf16.vhdl:300:40  */
  assign n1961 = x == 7'b1100000;
  /* fppowbf16.vhdl:301:40  */
  assign n1964 = x == 7'b1100001;
  /* fppowbf16.vhdl:302:40  */
  assign n1967 = x == 7'b1100010;
  /* fppowbf16.vhdl:303:40  */
  assign n1970 = x == 7'b1100011;
  /* fppowbf16.vhdl:304:40  */
  assign n1973 = x == 7'b1100100;
  /* fppowbf16.vhdl:305:40  */
  assign n1976 = x == 7'b1100101;
  /* fppowbf16.vhdl:306:40  */
  assign n1979 = x == 7'b1100110;
  /* fppowbf16.vhdl:307:40  */
  assign n1982 = x == 7'b1100111;
  /* fppowbf16.vhdl:308:40  */
  assign n1985 = x == 7'b1101000;
  /* fppowbf16.vhdl:309:40  */
  assign n1988 = x == 7'b1101001;
  /* fppowbf16.vhdl:310:40  */
  assign n1991 = x == 7'b1101010;
  /* fppowbf16.vhdl:311:40  */
  assign n1994 = x == 7'b1101011;
  /* fppowbf16.vhdl:312:40  */
  assign n1997 = x == 7'b1101100;
  /* fppowbf16.vhdl:313:40  */
  assign n2000 = x == 7'b1101101;
  /* fppowbf16.vhdl:314:40  */
  assign n2003 = x == 7'b1101110;
  /* fppowbf16.vhdl:315:40  */
  assign n2006 = x == 7'b1101111;
  /* fppowbf16.vhdl:316:40  */
  assign n2009 = x == 7'b1110000;
  /* fppowbf16.vhdl:317:40  */
  assign n2012 = x == 7'b1110001;
  /* fppowbf16.vhdl:318:40  */
  assign n2015 = x == 7'b1110010;
  /* fppowbf16.vhdl:319:40  */
  assign n2018 = x == 7'b1110011;
  /* fppowbf16.vhdl:320:40  */
  assign n2021 = x == 7'b1110100;
  /* fppowbf16.vhdl:321:40  */
  assign n2024 = x == 7'b1110101;
  /* fppowbf16.vhdl:322:40  */
  assign n2027 = x == 7'b1110110;
  /* fppowbf16.vhdl:323:40  */
  assign n2030 = x == 7'b1110111;
  /* fppowbf16.vhdl:324:40  */
  assign n2033 = x == 7'b1111000;
  /* fppowbf16.vhdl:325:40  */
  assign n2036 = x == 7'b1111001;
  /* fppowbf16.vhdl:326:40  */
  assign n2039 = x == 7'b1111010;
  /* fppowbf16.vhdl:327:40  */
  assign n2042 = x == 7'b1111011;
  /* fppowbf16.vhdl:328:40  */
  assign n2045 = x == 7'b1111100;
  /* fppowbf16.vhdl:329:40  */
  assign n2048 = x == 7'b1111101;
  /* fppowbf16.vhdl:330:40  */
  assign n2051 = x == 7'b1111110;
  /* fppowbf16.vhdl:331:40  */
  assign n2054 = x == 7'b1111111;
  assign n2056 = {n2054, n2051, n2048, n2045, n2042, n2039, n2036, n2033, n2030, n2027, n2024, n2021, n2018, n2015, n2012, n2009, n2006, n2003, n2000, n1997, n1994, n1991, n1988, n1985, n1982, n1979, n1976, n1973, n1970, n1967, n1964, n1961, n1958, n1955, n1952, n1949, n1946, n1943, n1940, n1937, n1934, n1931, n1928, n1925, n1922, n1919, n1916, n1913, n1910, n1907, n1904, n1901, n1898, n1895, n1892, n1889, n1886, n1883, n1880, n1877, n1874, n1871, n1868, n1865, n1862, n1859, n1856, n1853, n1850, n1847, n1844, n1841, n1838, n1835, n1832, n1829, n1826, n1823, n1820, n1817, n1814, n1811, n1808, n1805, n1802, n1799, n1796, n1793, n1790, n1787, n1784, n1781, n1778, n1775, n1772, n1769, n1766, n1763, n1760, n1757, n1754, n1751, n1748, n1745, n1742, n1739, n1736, n1733, n1730, n1727, n1724, n1721, n1718, n1715, n1712, n1709, n1706, n1703, n1700, n1697, n1694, n1691, n1688, n1685, n1682, n1679, n1676, n1673};
  /* fppowbf16.vhdl:203:4  */
  always @*
    case (n2056)
      128'b10000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2057 = 30'b111111011100000111111101010110;
      128'b01000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2057 = 30'b111110111100011111101010111010;
      128'b00100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2057 = 30'b111110111100011111101010111010;
      128'b00010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2057 = 30'b111110011101000110111001010000;
      128'b00001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2057 = 30'b111110011101000110111001010000;
      128'b00000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2057 = 30'b111101111101111101011001001111;
      128'b00000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2057 = 30'b111101111101111101011001001111;
      128'b00000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2057 = 30'b111101011111000010111100001001;
      128'b00000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2057 = 30'b111101011111000010111100001001;
      128'b00000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2057 = 30'b111101000000010111010011100001;
      128'b00000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2057 = 30'b111101000000010111010011100001;
      128'b00000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2057 = 30'b111100100001111010010001010010;
      128'b00000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2057 = 30'b111100100001111010010001010010;
      128'b00000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2057 = 30'b111100000011101011100111101000;
      128'b00000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2057 = 30'b111100000011101011100111101000;
      128'b00000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2057 = 30'b111011100101101011001001000100;
      128'b00000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2057 = 30'b111011000111111000101000011010;
      128'b00000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2057 = 30'b111011000111111000101000011010;
      128'b00000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2057 = 30'b111010101010010011111000110000;
      128'b00000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2057 = 30'b111010101010010011111000110000;
      128'b00000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2057 = 30'b111010001100111100101101011101;
      128'b00000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2057 = 30'b111001101111110010111010001010;
      128'b00000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2057 = 30'b111001101111110010111010001010;
      128'b00000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2057 = 30'b111001010010110110010010110001;
      128'b00000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2057 = 30'b111001010010110110010010110001;
      128'b00000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2057 = 30'b111000110110000110101011011100;
      128'b00000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2057 = 30'b111000011001100011111000100100;
      128'b00000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2057 = 30'b111000011001100011111000100100;
      128'b00000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2057 = 30'b110111111101001101101110110100;
      128'b00000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2057 = 30'b110111111101001101101110110100;
      128'b00000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2057 = 30'b110111100001000100000011000010;
      128'b00000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2057 = 30'b110111000101000110101010010110;
      128'b00000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2057 = 30'b110111000101000110101010010110;
      128'b00000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2057 = 30'b110110101001010101011010000100;
      128'b00000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2057 = 30'b110110001101110000000111110000;
      128'b00000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2057 = 30'b110110001101110000000111110000;
      128'b00000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2057 = 30'b110101110010010110101001001010;
      128'b00000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2057 = 30'b110101010111001000110100001110;
      128'b00000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2057 = 30'b110100111100000110011111001000;
      128'b00000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2057 = 30'b110100111100000110011111001000;
      128'b00000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2057 = 30'b110100100001001111100000001100;
      128'b00000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2057 = 30'b110100000110100011101101111111;
      128'b00000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2057 = 30'b110100000110100011101101111111;
      128'b00000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2057 = 30'b110011101100000010111111001110;
      128'b00000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2057 = 30'b110011010001101101001010110010;
      128'b00000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2057 = 30'b110010110111100010000111110000;
      128'b00000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2057 = 30'b110010110111100010000111110000;
      128'b00000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000: n2057 = 30'b110010011101100001101101011001;
      128'b00000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000: n2057 = 30'b110010000011101011110011000110;
      128'b00000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000: n2057 = 30'b110001101010000000010000011100;
      128'b00000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000: n2057 = 30'b110001101010000000010000011100;
      128'b00000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000: n2057 = 30'b110001010000011110111101001010;
      128'b00000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000: n2057 = 30'b110000110111000111110001001001;
      128'b00000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000: n2057 = 30'b110000011101111010100100011010;
      128'b00000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000: n2057 = 30'b110000000100110111001111001001;
      128'b00000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000: n2057 = 30'b110000000100110111001111001001;
      128'b00000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000: n2057 = 30'b101111101011111101101001101100;
      128'b00000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000: n2057 = 30'b101111010011001101101100011110;
      128'b00000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000: n2057 = 30'b101110111010100111010000000110;
      128'b00000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000: n2057 = 30'b101110100010001010001101010100;
      128'b00000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000: n2057 = 30'b101110001001110110011100111110;
      128'b00000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000: n2057 = 30'b101110001001110110011100111110;
      128'b00000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000: n2057 = 30'b101101110001101011111000000100;
      128'b00000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000: n2057 = 30'b101101011001101010010111101100;
      128'b00000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000: n2057 = 30'b011001011000111010001101000011;
      128'b00000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000: n2057 = 30'b011000101001100011100110101000;
      128'b00000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000: n2057 = 30'b011000101001100011100110101000;
      128'b00000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000: n2057 = 30'b010111111010101111101000111100;
      128'b00000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000: n2057 = 30'b010111111010101111101000111100;
      128'b00000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000: n2057 = 30'b010111001100011101100001110111;
      128'b00000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000: n2057 = 30'b010111001100011101100001110111;
      128'b00000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000: n2057 = 30'b010110011110101100100000111110;
      128'b00000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000: n2057 = 30'b010110011110101100100000111110;
      128'b00000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000: n2057 = 30'b010101110001011011110111100000;
      128'b00000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000: n2057 = 30'b010101110001011011110111100000;
      128'b00000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000: n2057 = 30'b010101000100101010111000000111;
      128'b00000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000: n2057 = 30'b010101000100101010111000000111;
      128'b00000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000: n2057 = 30'b010100011000011000110111000010;
      128'b00000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000: n2057 = 30'b010100011000011000110111000010;
      128'b00000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000: n2057 = 30'b010011101100100101001001110111;
      128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000: n2057 = 30'b010011101100100101001001110111;
      128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000: n2057 = 30'b010011000001001111000111100010;
      128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000: n2057 = 30'b010011000001001111000111100010;
      128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000: n2057 = 30'b010010010110010110001000010001;
      128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000: n2057 = 30'b010010010110010110001000010001;
      128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000: n2057 = 30'b010001101011111001100101100100;
      128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000: n2057 = 30'b010001101011111001100101100100;
      128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000: n2057 = 30'b010001000001111000111010000010;
      128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000: n2057 = 30'b010000011000010011100001100000;
      128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000: n2057 = 30'b010000011000010011100001100000;
      128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000: n2057 = 30'b001111101111001000111000110110;
      128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000: n2057 = 30'b001111101111001000111000110110;
      128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000: n2057 = 30'b001111000110011000011110000000;
      128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000: n2057 = 30'b001110011110000001101111111001;
      128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000: n2057 = 30'b001110011110000001101111111001;
      128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000: n2057 = 30'b001101110110000100001110011100;
      128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000: n2057 = 30'b001101001110011111011010011110;
      128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000: n2057 = 30'b001101001110011111011010011110;
      128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000: n2057 = 30'b001100100111010010110101101110;
      128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000: n2057 = 30'b001100000000011110000010110011;
      128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000: n2057 = 30'b001100000000011110000010110011;
      128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000: n2057 = 30'b001011011010000000100101000110;
      128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000: n2057 = 30'b001010110011111010000000110110;
      128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000: n2057 = 30'b001010110011111010000000110110;
      128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000: n2057 = 30'b001010001110001001111011000010;
      128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000: n2057 = 30'b001001101000101111111001011000;
      128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000: n2057 = 30'b001001101000101111111001011000;
      128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000: n2057 = 30'b001001000011101011100010010101;
      128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000: n2057 = 30'b001000011110111100011101000001;
      128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000: n2057 = 30'b000111111010100010010001001110;
      128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000: n2057 = 30'b000111111010100010010001001110;
      128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000: n2057 = 30'b000111010110011100100111011001;
      128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000: n2057 = 30'b000110110010101011001000100011;
      128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000: n2057 = 30'b000110001111001101011110010111;
      128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000: n2057 = 30'b000101101100000011010011000011;
      128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000: n2057 = 30'b000101001001001100010001010111;
      128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000: n2057 = 30'b000101001001001100010001010111;
      128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000: n2057 = 30'b000100100110101000000100101001;
      128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000: n2057 = 30'b000100000100010110011000101101;
      128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000: n2057 = 30'b000011100010010110111001111010;
      128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000: n2057 = 30'b000011000000101001010101000011;
      128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000: n2057 = 30'b000010011111001101010111011010;
      128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000: n2057 = 30'b000001111110000010101110110001;
      128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000: n2057 = 30'b000001011101001001001001010011;
      128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000: n2057 = 30'b000000111100100000010101100110;
      128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100: n2057 = 30'b000000011100001000000010101100;
      128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010: n2057 = 30'b111111111100000000000000000000;
      128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001: n2057 = 30'b111111111100000000000000000000;
      default: n2057 = 30'bX;
    endcase
endmodule

module intadder_21_freq500_uid25
  (input  clk,
   input  [20:0] x,
   input  [20:0] y,
   input  cin,
   output [20:0] r);
  wire [20:0] rtmp;
  wire [20:0] x_d1;
  wire [20:0] x_d2;
  wire [20:0] x_d3;
  wire [20:0] y_d1;
  wire cin_d1;
  wire cin_d2;
  wire cin_d3;
  wire cin_d4;
  wire cin_d5;
  wire cin_d6;
  wire [20:0] n1657;
  wire [20:0] n1658;
  wire [20:0] n1659;
  reg [20:0] n1660;
  reg [20:0] n1661;
  reg [20:0] n1662;
  reg [20:0] n1663;
  reg n1664;
  reg n1665;
  reg n1666;
  reg n1667;
  reg n1668;
  reg n1669;
  assign r = rtmp; //(module output)
  /* fppowbf16.vhdl:2266:8  */
  assign rtmp = n1659; // (signal)
  /* fppowbf16.vhdl:2268:8  */
  assign x_d1 = n1660; // (signal)
  /* fppowbf16.vhdl:2268:14  */
  assign x_d2 = n1661; // (signal)
  /* fppowbf16.vhdl:2268:20  */
  assign x_d3 = n1662; // (signal)
  /* fppowbf16.vhdl:2270:8  */
  assign y_d1 = n1663; // (signal)
  /* fppowbf16.vhdl:2272:8  */
  assign cin_d1 = n1664; // (signal)
  /* fppowbf16.vhdl:2272:16  */
  assign cin_d2 = n1665; // (signal)
  /* fppowbf16.vhdl:2272:24  */
  assign cin_d3 = n1666; // (signal)
  /* fppowbf16.vhdl:2272:32  */
  assign cin_d4 = n1667; // (signal)
  /* fppowbf16.vhdl:2272:40  */
  assign cin_d5 = n1668; // (signal)
  /* fppowbf16.vhdl:2272:48  */
  assign cin_d6 = n1669; // (signal)
  /* fppowbf16.vhdl:2290:17  */
  assign n1657 = x_d3 + y_d1;
  /* fppowbf16.vhdl:2290:24  */
  assign n1658 = {20'b0, cin_d6};  //  uext
  /* fppowbf16.vhdl:2290:24  */
  assign n1659 = n1657 + n1658;
  /* fppowbf16.vhdl:2277:10  */
  always @(posedge clk)
    n1660 <= x;
  /* fppowbf16.vhdl:2277:10  */
  always @(posedge clk)
    n1661 <= x_d1;
  /* fppowbf16.vhdl:2277:10  */
  always @(posedge clk)
    n1662 <= x_d2;
  /* fppowbf16.vhdl:2277:10  */
  always @(posedge clk)
    n1663 <= y;
  /* fppowbf16.vhdl:2277:10  */
  always @(posedge clk)
    n1664 <= cin;
  /* fppowbf16.vhdl:2277:10  */
  always @(posedge clk)
    n1665 <= cin_d1;
  /* fppowbf16.vhdl:2277:10  */
  always @(posedge clk)
    n1666 <= cin_d2;
  /* fppowbf16.vhdl:2277:10  */
  always @(posedge clk)
    n1667 <= cin_d3;
  /* fppowbf16.vhdl:2277:10  */
  always @(posedge clk)
    n1668 <= cin_d4;
  /* fppowbf16.vhdl:2277:10  */
  always @(posedge clk)
    n1669 <= cin_d5;
endmodule

module intadder_21_freq500_uid22
  (input  clk,
   input  [20:0] x,
   input  [20:0] y,
   input  cin,
   output [20:0] r);
  wire cin_1;
  wire cin_1_d1;
  wire cin_1_d2;
  wire cin_1_d3;
  wire [21:0] x_1;
  wire [21:0] x_1_d1;
  wire [21:0] y_1;
  wire [21:0] y_1_d1;
  wire [21:0] s_1;
  wire [20:0] r_1;
  wire [21:0] n1630;
  wire [21:0] n1632;
  wire [21:0] n1633;
  wire [21:0] n1634;
  wire [21:0] n1635;
  wire [20:0] n1636;
  reg n1637;
  reg n1638;
  reg n1639;
  reg [21:0] n1640;
  reg [21:0] n1641;
  assign r = r_1; //(module output)
  /* fppowbf16.vhdl:2205:15  */
  assign cin_1_d1 = n1637; // (signal)
  /* fppowbf16.vhdl:2205:25  */
  assign cin_1_d2 = n1638; // (signal)
  /* fppowbf16.vhdl:2205:35  */
  assign cin_1_d3 = n1639; // (signal)
  /* fppowbf16.vhdl:2207:8  */
  assign x_1 = n1630; // (signal)
  /* fppowbf16.vhdl:2207:13  */
  assign x_1_d1 = n1640; // (signal)
  /* fppowbf16.vhdl:2209:8  */
  assign y_1 = n1632; // (signal)
  /* fppowbf16.vhdl:2209:13  */
  assign y_1_d1 = n1641; // (signal)
  /* fppowbf16.vhdl:2211:8  */
  assign s_1 = n1635; // (signal)
  /* fppowbf16.vhdl:2213:8  */
  assign r_1 = n1636; // (signal)
  /* fppowbf16.vhdl:2227:15  */
  assign n1630 = {1'b0, x};
  /* fppowbf16.vhdl:2228:15  */
  assign n1632 = {1'b0, y};
  /* fppowbf16.vhdl:2229:18  */
  assign n1633 = x_1_d1 + y_1_d1;
  /* fppowbf16.vhdl:2229:27  */
  assign n1634 = {21'b0, cin_1_d3};  //  uext
  /* fppowbf16.vhdl:2229:27  */
  assign n1635 = n1633 + n1634;
  /* fppowbf16.vhdl:2230:14  */
  assign n1636 = s_1[20:0]; // extract
  /* fppowbf16.vhdl:2218:10  */
  always @(posedge clk)
    n1637 <= cin_1;
  /* fppowbf16.vhdl:2218:10  */
  always @(posedge clk)
    n1638 <= cin_1_d1;
  /* fppowbf16.vhdl:2218:10  */
  always @(posedge clk)
    n1639 <= cin_1_d2;
  /* fppowbf16.vhdl:2218:10  */
  always @(posedge clk)
    n1640 <= x_1;
  /* fppowbf16.vhdl:2218:10  */
  always @(posedge clk)
    n1641 <= y_1;
endmodule

module intadder_21_freq500_uid19
  (input  clk,
   input  [20:0] x,
   input  [20:0] y,
   input  cin,
   output [20:0] r);
  wire cin_1;
  wire cin_1_d1;
  wire cin_1_d2;
  wire [21:0] x_1;
  wire [21:0] x_1_d1;
  wire [21:0] y_1;
  wire [21:0] y_1_d1;
  wire [21:0] s_1;
  wire [20:0] r_1;
  wire [21:0] n1608;
  wire [21:0] n1610;
  wire [21:0] n1611;
  wire [21:0] n1612;
  wire [21:0] n1613;
  wire [20:0] n1614;
  reg n1615;
  reg n1616;
  reg [21:0] n1617;
  reg [21:0] n1618;
  assign r = r_1; //(module output)
  /* fppowbf16.vhdl:2145:15  */
  assign cin_1_d1 = n1615; // (signal)
  /* fppowbf16.vhdl:2145:25  */
  assign cin_1_d2 = n1616; // (signal)
  /* fppowbf16.vhdl:2147:8  */
  assign x_1 = n1608; // (signal)
  /* fppowbf16.vhdl:2147:13  */
  assign x_1_d1 = n1617; // (signal)
  /* fppowbf16.vhdl:2149:8  */
  assign y_1 = n1610; // (signal)
  /* fppowbf16.vhdl:2149:13  */
  assign y_1_d1 = n1618; // (signal)
  /* fppowbf16.vhdl:2151:8  */
  assign s_1 = n1613; // (signal)
  /* fppowbf16.vhdl:2153:8  */
  assign r_1 = n1614; // (signal)
  /* fppowbf16.vhdl:2166:15  */
  assign n1608 = {1'b0, x};
  /* fppowbf16.vhdl:2167:15  */
  assign n1610 = {1'b0, y};
  /* fppowbf16.vhdl:2168:18  */
  assign n1611 = x_1_d1 + y_1_d1;
  /* fppowbf16.vhdl:2168:27  */
  assign n1612 = {21'b0, cin_1_d2};  //  uext
  /* fppowbf16.vhdl:2168:27  */
  assign n1613 = n1611 + n1612;
  /* fppowbf16.vhdl:2169:14  */
  assign n1614 = s_1[20:0]; // extract
  /* fppowbf16.vhdl:2158:10  */
  always @(posedge clk)
    n1615 <= cin_1;
  /* fppowbf16.vhdl:2158:10  */
  always @(posedge clk)
    n1616 <= cin_1_d1;
  /* fppowbf16.vhdl:2158:10  */
  always @(posedge clk)
    n1617 <= x_1;
  /* fppowbf16.vhdl:2158:10  */
  always @(posedge clk)
    n1618 <= y_1;
endmodule

module inva0table_freq500_uid15
  (input  [6:0] x,
   output [7:0] y);
  wire [7:0] y0;
  wire [7:0] y1;
  wire n1213;
  wire n1216;
  wire n1219;
  wire n1222;
  wire n1225;
  wire n1228;
  wire n1231;
  wire n1234;
  wire n1237;
  wire n1240;
  wire n1243;
  wire n1246;
  wire n1249;
  wire n1252;
  wire n1255;
  wire n1258;
  wire n1261;
  wire n1264;
  wire n1267;
  wire n1270;
  wire n1273;
  wire n1276;
  wire n1279;
  wire n1282;
  wire n1285;
  wire n1288;
  wire n1291;
  wire n1294;
  wire n1297;
  wire n1300;
  wire n1303;
  wire n1306;
  wire n1309;
  wire n1312;
  wire n1315;
  wire n1318;
  wire n1321;
  wire n1324;
  wire n1327;
  wire n1330;
  wire n1333;
  wire n1336;
  wire n1339;
  wire n1342;
  wire n1345;
  wire n1348;
  wire n1351;
  wire n1354;
  wire n1357;
  wire n1360;
  wire n1363;
  wire n1366;
  wire n1369;
  wire n1372;
  wire n1375;
  wire n1378;
  wire n1381;
  wire n1384;
  wire n1387;
  wire n1390;
  wire n1393;
  wire n1396;
  wire n1399;
  wire n1402;
  wire n1405;
  wire n1408;
  wire n1411;
  wire n1414;
  wire n1417;
  wire n1420;
  wire n1423;
  wire n1426;
  wire n1429;
  wire n1432;
  wire n1435;
  wire n1438;
  wire n1441;
  wire n1444;
  wire n1447;
  wire n1450;
  wire n1453;
  wire n1456;
  wire n1459;
  wire n1462;
  wire n1465;
  wire n1468;
  wire n1471;
  wire n1474;
  wire n1477;
  wire n1480;
  wire n1483;
  wire n1486;
  wire n1489;
  wire n1492;
  wire n1495;
  wire n1498;
  wire n1501;
  wire n1504;
  wire n1507;
  wire n1510;
  wire n1513;
  wire n1516;
  wire n1519;
  wire n1522;
  wire n1525;
  wire n1528;
  wire n1531;
  wire n1534;
  wire n1537;
  wire n1540;
  wire n1543;
  wire n1546;
  wire n1549;
  wire n1552;
  wire n1555;
  wire n1558;
  wire n1561;
  wire n1564;
  wire n1567;
  wire n1570;
  wire n1573;
  wire n1576;
  wire n1579;
  wire n1582;
  wire n1585;
  wire n1588;
  wire n1591;
  wire n1594;
  wire [127:0] n1596;
  reg [7:0] n1597;
  assign y = y1; //(module output)
  /* fppowbf16.vhdl:30:8  */
  assign y0 = n1597; // (signal)
  /* fppowbf16.vhdl:32:8  */
  assign y1 = y0; // (signal)
  /* fppowbf16.vhdl:36:18  */
  assign n1213 = x == 7'b0000000;
  /* fppowbf16.vhdl:37:18  */
  assign n1216 = x == 7'b0000001;
  /* fppowbf16.vhdl:38:18  */
  assign n1219 = x == 7'b0000010;
  /* fppowbf16.vhdl:39:18  */
  assign n1222 = x == 7'b0000011;
  /* fppowbf16.vhdl:40:18  */
  assign n1225 = x == 7'b0000100;
  /* fppowbf16.vhdl:41:18  */
  assign n1228 = x == 7'b0000101;
  /* fppowbf16.vhdl:42:18  */
  assign n1231 = x == 7'b0000110;
  /* fppowbf16.vhdl:43:18  */
  assign n1234 = x == 7'b0000111;
  /* fppowbf16.vhdl:44:18  */
  assign n1237 = x == 7'b0001000;
  /* fppowbf16.vhdl:45:18  */
  assign n1240 = x == 7'b0001001;
  /* fppowbf16.vhdl:46:18  */
  assign n1243 = x == 7'b0001010;
  /* fppowbf16.vhdl:47:18  */
  assign n1246 = x == 7'b0001011;
  /* fppowbf16.vhdl:48:18  */
  assign n1249 = x == 7'b0001100;
  /* fppowbf16.vhdl:49:18  */
  assign n1252 = x == 7'b0001101;
  /* fppowbf16.vhdl:50:18  */
  assign n1255 = x == 7'b0001110;
  /* fppowbf16.vhdl:51:18  */
  assign n1258 = x == 7'b0001111;
  /* fppowbf16.vhdl:52:18  */
  assign n1261 = x == 7'b0010000;
  /* fppowbf16.vhdl:53:18  */
  assign n1264 = x == 7'b0010001;
  /* fppowbf16.vhdl:54:18  */
  assign n1267 = x == 7'b0010010;
  /* fppowbf16.vhdl:55:18  */
  assign n1270 = x == 7'b0010011;
  /* fppowbf16.vhdl:56:18  */
  assign n1273 = x == 7'b0010100;
  /* fppowbf16.vhdl:57:18  */
  assign n1276 = x == 7'b0010101;
  /* fppowbf16.vhdl:58:18  */
  assign n1279 = x == 7'b0010110;
  /* fppowbf16.vhdl:59:18  */
  assign n1282 = x == 7'b0010111;
  /* fppowbf16.vhdl:60:18  */
  assign n1285 = x == 7'b0011000;
  /* fppowbf16.vhdl:61:18  */
  assign n1288 = x == 7'b0011001;
  /* fppowbf16.vhdl:62:18  */
  assign n1291 = x == 7'b0011010;
  /* fppowbf16.vhdl:63:18  */
  assign n1294 = x == 7'b0011011;
  /* fppowbf16.vhdl:64:18  */
  assign n1297 = x == 7'b0011100;
  /* fppowbf16.vhdl:65:18  */
  assign n1300 = x == 7'b0011101;
  /* fppowbf16.vhdl:66:18  */
  assign n1303 = x == 7'b0011110;
  /* fppowbf16.vhdl:67:18  */
  assign n1306 = x == 7'b0011111;
  /* fppowbf16.vhdl:68:18  */
  assign n1309 = x == 7'b0100000;
  /* fppowbf16.vhdl:69:18  */
  assign n1312 = x == 7'b0100001;
  /* fppowbf16.vhdl:70:18  */
  assign n1315 = x == 7'b0100010;
  /* fppowbf16.vhdl:71:18  */
  assign n1318 = x == 7'b0100011;
  /* fppowbf16.vhdl:72:18  */
  assign n1321 = x == 7'b0100100;
  /* fppowbf16.vhdl:73:18  */
  assign n1324 = x == 7'b0100101;
  /* fppowbf16.vhdl:74:18  */
  assign n1327 = x == 7'b0100110;
  /* fppowbf16.vhdl:75:18  */
  assign n1330 = x == 7'b0100111;
  /* fppowbf16.vhdl:76:18  */
  assign n1333 = x == 7'b0101000;
  /* fppowbf16.vhdl:77:18  */
  assign n1336 = x == 7'b0101001;
  /* fppowbf16.vhdl:78:18  */
  assign n1339 = x == 7'b0101010;
  /* fppowbf16.vhdl:79:18  */
  assign n1342 = x == 7'b0101011;
  /* fppowbf16.vhdl:80:18  */
  assign n1345 = x == 7'b0101100;
  /* fppowbf16.vhdl:81:18  */
  assign n1348 = x == 7'b0101101;
  /* fppowbf16.vhdl:82:18  */
  assign n1351 = x == 7'b0101110;
  /* fppowbf16.vhdl:83:18  */
  assign n1354 = x == 7'b0101111;
  /* fppowbf16.vhdl:84:18  */
  assign n1357 = x == 7'b0110000;
  /* fppowbf16.vhdl:85:18  */
  assign n1360 = x == 7'b0110001;
  /* fppowbf16.vhdl:86:18  */
  assign n1363 = x == 7'b0110010;
  /* fppowbf16.vhdl:87:18  */
  assign n1366 = x == 7'b0110011;
  /* fppowbf16.vhdl:88:18  */
  assign n1369 = x == 7'b0110100;
  /* fppowbf16.vhdl:89:18  */
  assign n1372 = x == 7'b0110101;
  /* fppowbf16.vhdl:90:18  */
  assign n1375 = x == 7'b0110110;
  /* fppowbf16.vhdl:91:18  */
  assign n1378 = x == 7'b0110111;
  /* fppowbf16.vhdl:92:18  */
  assign n1381 = x == 7'b0111000;
  /* fppowbf16.vhdl:93:18  */
  assign n1384 = x == 7'b0111001;
  /* fppowbf16.vhdl:94:18  */
  assign n1387 = x == 7'b0111010;
  /* fppowbf16.vhdl:95:18  */
  assign n1390 = x == 7'b0111011;
  /* fppowbf16.vhdl:96:18  */
  assign n1393 = x == 7'b0111100;
  /* fppowbf16.vhdl:97:18  */
  assign n1396 = x == 7'b0111101;
  /* fppowbf16.vhdl:98:18  */
  assign n1399 = x == 7'b0111110;
  /* fppowbf16.vhdl:99:18  */
  assign n1402 = x == 7'b0111111;
  /* fppowbf16.vhdl:100:18  */
  assign n1405 = x == 7'b1000000;
  /* fppowbf16.vhdl:101:18  */
  assign n1408 = x == 7'b1000001;
  /* fppowbf16.vhdl:102:18  */
  assign n1411 = x == 7'b1000010;
  /* fppowbf16.vhdl:103:18  */
  assign n1414 = x == 7'b1000011;
  /* fppowbf16.vhdl:104:18  */
  assign n1417 = x == 7'b1000100;
  /* fppowbf16.vhdl:105:18  */
  assign n1420 = x == 7'b1000101;
  /* fppowbf16.vhdl:106:18  */
  assign n1423 = x == 7'b1000110;
  /* fppowbf16.vhdl:107:18  */
  assign n1426 = x == 7'b1000111;
  /* fppowbf16.vhdl:108:18  */
  assign n1429 = x == 7'b1001000;
  /* fppowbf16.vhdl:109:18  */
  assign n1432 = x == 7'b1001001;
  /* fppowbf16.vhdl:110:18  */
  assign n1435 = x == 7'b1001010;
  /* fppowbf16.vhdl:111:18  */
  assign n1438 = x == 7'b1001011;
  /* fppowbf16.vhdl:112:18  */
  assign n1441 = x == 7'b1001100;
  /* fppowbf16.vhdl:113:18  */
  assign n1444 = x == 7'b1001101;
  /* fppowbf16.vhdl:114:18  */
  assign n1447 = x == 7'b1001110;
  /* fppowbf16.vhdl:115:18  */
  assign n1450 = x == 7'b1001111;
  /* fppowbf16.vhdl:116:18  */
  assign n1453 = x == 7'b1010000;
  /* fppowbf16.vhdl:117:18  */
  assign n1456 = x == 7'b1010001;
  /* fppowbf16.vhdl:118:18  */
  assign n1459 = x == 7'b1010010;
  /* fppowbf16.vhdl:119:18  */
  assign n1462 = x == 7'b1010011;
  /* fppowbf16.vhdl:120:18  */
  assign n1465 = x == 7'b1010100;
  /* fppowbf16.vhdl:121:18  */
  assign n1468 = x == 7'b1010101;
  /* fppowbf16.vhdl:122:18  */
  assign n1471 = x == 7'b1010110;
  /* fppowbf16.vhdl:123:18  */
  assign n1474 = x == 7'b1010111;
  /* fppowbf16.vhdl:124:18  */
  assign n1477 = x == 7'b1011000;
  /* fppowbf16.vhdl:125:18  */
  assign n1480 = x == 7'b1011001;
  /* fppowbf16.vhdl:126:18  */
  assign n1483 = x == 7'b1011010;
  /* fppowbf16.vhdl:127:18  */
  assign n1486 = x == 7'b1011011;
  /* fppowbf16.vhdl:128:18  */
  assign n1489 = x == 7'b1011100;
  /* fppowbf16.vhdl:129:18  */
  assign n1492 = x == 7'b1011101;
  /* fppowbf16.vhdl:130:18  */
  assign n1495 = x == 7'b1011110;
  /* fppowbf16.vhdl:131:18  */
  assign n1498 = x == 7'b1011111;
  /* fppowbf16.vhdl:132:18  */
  assign n1501 = x == 7'b1100000;
  /* fppowbf16.vhdl:133:18  */
  assign n1504 = x == 7'b1100001;
  /* fppowbf16.vhdl:134:18  */
  assign n1507 = x == 7'b1100010;
  /* fppowbf16.vhdl:135:18  */
  assign n1510 = x == 7'b1100011;
  /* fppowbf16.vhdl:136:18  */
  assign n1513 = x == 7'b1100100;
  /* fppowbf16.vhdl:137:18  */
  assign n1516 = x == 7'b1100101;
  /* fppowbf16.vhdl:138:18  */
  assign n1519 = x == 7'b1100110;
  /* fppowbf16.vhdl:139:18  */
  assign n1522 = x == 7'b1100111;
  /* fppowbf16.vhdl:140:18  */
  assign n1525 = x == 7'b1101000;
  /* fppowbf16.vhdl:141:18  */
  assign n1528 = x == 7'b1101001;
  /* fppowbf16.vhdl:142:18  */
  assign n1531 = x == 7'b1101010;
  /* fppowbf16.vhdl:143:18  */
  assign n1534 = x == 7'b1101011;
  /* fppowbf16.vhdl:144:18  */
  assign n1537 = x == 7'b1101100;
  /* fppowbf16.vhdl:145:18  */
  assign n1540 = x == 7'b1101101;
  /* fppowbf16.vhdl:146:18  */
  assign n1543 = x == 7'b1101110;
  /* fppowbf16.vhdl:147:18  */
  assign n1546 = x == 7'b1101111;
  /* fppowbf16.vhdl:148:18  */
  assign n1549 = x == 7'b1110000;
  /* fppowbf16.vhdl:149:18  */
  assign n1552 = x == 7'b1110001;
  /* fppowbf16.vhdl:150:18  */
  assign n1555 = x == 7'b1110010;
  /* fppowbf16.vhdl:151:18  */
  assign n1558 = x == 7'b1110011;
  /* fppowbf16.vhdl:152:18  */
  assign n1561 = x == 7'b1110100;
  /* fppowbf16.vhdl:153:18  */
  assign n1564 = x == 7'b1110101;
  /* fppowbf16.vhdl:154:18  */
  assign n1567 = x == 7'b1110110;
  /* fppowbf16.vhdl:155:18  */
  assign n1570 = x == 7'b1110111;
  /* fppowbf16.vhdl:156:18  */
  assign n1573 = x == 7'b1111000;
  /* fppowbf16.vhdl:157:18  */
  assign n1576 = x == 7'b1111001;
  /* fppowbf16.vhdl:158:18  */
  assign n1579 = x == 7'b1111010;
  /* fppowbf16.vhdl:159:18  */
  assign n1582 = x == 7'b1111011;
  /* fppowbf16.vhdl:160:18  */
  assign n1585 = x == 7'b1111100;
  /* fppowbf16.vhdl:161:18  */
  assign n1588 = x == 7'b1111101;
  /* fppowbf16.vhdl:162:18  */
  assign n1591 = x == 7'b1111110;
  /* fppowbf16.vhdl:163:18  */
  assign n1594 = x == 7'b1111111;
  assign n1596 = {n1594, n1591, n1588, n1585, n1582, n1579, n1576, n1573, n1570, n1567, n1564, n1561, n1558, n1555, n1552, n1549, n1546, n1543, n1540, n1537, n1534, n1531, n1528, n1525, n1522, n1519, n1516, n1513, n1510, n1507, n1504, n1501, n1498, n1495, n1492, n1489, n1486, n1483, n1480, n1477, n1474, n1471, n1468, n1465, n1462, n1459, n1456, n1453, n1450, n1447, n1444, n1441, n1438, n1435, n1432, n1429, n1426, n1423, n1420, n1417, n1414, n1411, n1408, n1405, n1402, n1399, n1396, n1393, n1390, n1387, n1384, n1381, n1378, n1375, n1372, n1369, n1366, n1363, n1360, n1357, n1354, n1351, n1348, n1345, n1342, n1339, n1336, n1333, n1330, n1327, n1324, n1321, n1318, n1315, n1312, n1309, n1306, n1303, n1300, n1297, n1294, n1291, n1288, n1285, n1282, n1279, n1276, n1273, n1270, n1267, n1264, n1261, n1258, n1255, n1252, n1249, n1246, n1243, n1240, n1237, n1234, n1231, n1228, n1225, n1222, n1219, n1216, n1213};
  /* fppowbf16.vhdl:35:4  */
  always @*
    case (n1596)
      128'b10000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1597 = 8'b10000001;
      128'b01000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1597 = 8'b10000010;
      128'b00100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1597 = 8'b10000010;
      128'b00010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1597 = 8'b10000011;
      128'b00001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1597 = 8'b10000011;
      128'b00000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1597 = 8'b10000100;
      128'b00000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1597 = 8'b10000100;
      128'b00000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1597 = 8'b10000101;
      128'b00000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1597 = 8'b10000101;
      128'b00000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1597 = 8'b10000110;
      128'b00000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1597 = 8'b10000110;
      128'b00000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1597 = 8'b10000111;
      128'b00000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1597 = 8'b10000111;
      128'b00000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1597 = 8'b10001000;
      128'b00000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1597 = 8'b10001000;
      128'b00000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1597 = 8'b10001001;
      128'b00000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1597 = 8'b10001010;
      128'b00000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1597 = 8'b10001010;
      128'b00000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1597 = 8'b10001011;
      128'b00000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1597 = 8'b10001011;
      128'b00000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1597 = 8'b10001100;
      128'b00000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1597 = 8'b10001101;
      128'b00000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1597 = 8'b10001101;
      128'b00000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1597 = 8'b10001110;
      128'b00000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1597 = 8'b10001110;
      128'b00000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1597 = 8'b10001111;
      128'b00000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1597 = 8'b10010000;
      128'b00000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1597 = 8'b10010000;
      128'b00000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1597 = 8'b10010001;
      128'b00000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1597 = 8'b10010001;
      128'b00000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1597 = 8'b10010010;
      128'b00000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1597 = 8'b10010011;
      128'b00000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1597 = 8'b10010011;
      128'b00000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1597 = 8'b10010100;
      128'b00000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1597 = 8'b10010101;
      128'b00000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1597 = 8'b10010101;
      128'b00000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1597 = 8'b10010110;
      128'b00000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1597 = 8'b10010111;
      128'b00000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1597 = 8'b10011000;
      128'b00000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1597 = 8'b10011000;
      128'b00000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1597 = 8'b10011001;
      128'b00000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1597 = 8'b10011010;
      128'b00000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1597 = 8'b10011010;
      128'b00000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1597 = 8'b10011011;
      128'b00000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1597 = 8'b10011100;
      128'b00000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1597 = 8'b10011101;
      128'b00000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1597 = 8'b10011101;
      128'b00000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000: n1597 = 8'b10011110;
      128'b00000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000: n1597 = 8'b10011111;
      128'b00000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000: n1597 = 8'b10100000;
      128'b00000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000: n1597 = 8'b10100000;
      128'b00000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000: n1597 = 8'b10100001;
      128'b00000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000: n1597 = 8'b10100010;
      128'b00000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000: n1597 = 8'b10100011;
      128'b00000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000: n1597 = 8'b10100100;
      128'b00000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000: n1597 = 8'b10100100;
      128'b00000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000: n1597 = 8'b10100101;
      128'b00000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000: n1597 = 8'b10100110;
      128'b00000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000: n1597 = 8'b10100111;
      128'b00000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000: n1597 = 8'b10101000;
      128'b00000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000: n1597 = 8'b10101001;
      128'b00000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000: n1597 = 8'b10101001;
      128'b00000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000: n1597 = 8'b10101010;
      128'b00000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000: n1597 = 8'b10101011;
      128'b00000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000: n1597 = 8'b01010110;
      128'b00000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000: n1597 = 8'b01010111;
      128'b00000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000: n1597 = 8'b01010111;
      128'b00000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000: n1597 = 8'b01011000;
      128'b00000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000: n1597 = 8'b01011000;
      128'b00000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000: n1597 = 8'b01011001;
      128'b00000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000: n1597 = 8'b01011001;
      128'b00000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000: n1597 = 8'b01011010;
      128'b00000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000: n1597 = 8'b01011010;
      128'b00000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000: n1597 = 8'b01011011;
      128'b00000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000: n1597 = 8'b01011011;
      128'b00000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000: n1597 = 8'b01011100;
      128'b00000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000: n1597 = 8'b01011100;
      128'b00000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000: n1597 = 8'b01011101;
      128'b00000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000: n1597 = 8'b01011101;
      128'b00000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000: n1597 = 8'b01011110;
      128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000: n1597 = 8'b01011110;
      128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000: n1597 = 8'b01011111;
      128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000: n1597 = 8'b01011111;
      128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000: n1597 = 8'b01100000;
      128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000: n1597 = 8'b01100000;
      128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000: n1597 = 8'b01100001;
      128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000: n1597 = 8'b01100001;
      128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000: n1597 = 8'b01100010;
      128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000: n1597 = 8'b01100011;
      128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000: n1597 = 8'b01100011;
      128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000: n1597 = 8'b01100100;
      128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000: n1597 = 8'b01100100;
      128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000: n1597 = 8'b01100101;
      128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000: n1597 = 8'b01100110;
      128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000: n1597 = 8'b01100110;
      128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000: n1597 = 8'b01100111;
      128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000: n1597 = 8'b01101000;
      128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000: n1597 = 8'b01101000;
      128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000: n1597 = 8'b01101001;
      128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000: n1597 = 8'b01101010;
      128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000: n1597 = 8'b01101010;
      128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000: n1597 = 8'b01101011;
      128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000: n1597 = 8'b01101100;
      128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000: n1597 = 8'b01101100;
      128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000: n1597 = 8'b01101101;
      128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000: n1597 = 8'b01101110;
      128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000: n1597 = 8'b01101110;
      128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000: n1597 = 8'b01101111;
      128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000: n1597 = 8'b01110000;
      128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000: n1597 = 8'b01110001;
      128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000: n1597 = 8'b01110001;
      128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000: n1597 = 8'b01110010;
      128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000: n1597 = 8'b01110011;
      128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000: n1597 = 8'b01110100;
      128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000: n1597 = 8'b01110101;
      128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000: n1597 = 8'b01110110;
      128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000: n1597 = 8'b01110110;
      128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000: n1597 = 8'b01110111;
      128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000: n1597 = 8'b01111000;
      128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000: n1597 = 8'b01111001;
      128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000: n1597 = 8'b01111010;
      128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000: n1597 = 8'b01111011;
      128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000: n1597 = 8'b01111100;
      128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000: n1597 = 8'b01111101;
      128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000: n1597 = 8'b01111110;
      128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100: n1597 = 8'b01111111;
      128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010: n1597 = 8'b10000000;
      128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001: n1597 = 8'b10000000;
      default: n1597 = 8'bX;
    endcase
endmodule

module leftshifter10_by_max_10_freq500_uid13
  (input  clk,
   input  [9:0] x,
   input  [3:0] s,
   output [19:0] r);
  wire [3:0] ps;
  wire [3:0] ps_d1;
  wire [9:0] level0;
  wire [9:0] level0_d1;
  wire [9:0] level0_d2;
  wire [9:0] level0_d3;
  wire [10:0] level1;
  wire [10:0] level1_d1;
  wire [12:0] level2;
  wire [16:0] level3;
  wire [24:0] level4;
  wire [10:0] n1181;
  wire n1182;
  wire [10:0] n1183;
  wire [10:0] n1185;
  wire [12:0] n1187;
  wire n1188;
  wire [12:0] n1189;
  wire [12:0] n1191;
  wire [16:0] n1193;
  wire n1194;
  wire [16:0] n1195;
  wire [16:0] n1197;
  wire [24:0] n1199;
  wire n1200;
  wire [24:0] n1201;
  wire [24:0] n1203;
  wire [19:0] n1204;
  reg [3:0] n1205;
  reg [9:0] n1206;
  reg [9:0] n1207;
  reg [9:0] n1208;
  reg [10:0] n1209;
  assign r = n1204; //(module output)
  /* fppowbf16.vhdl:2081:12  */
  assign ps_d1 = n1205; // (signal)
  /* fppowbf16.vhdl:2083:16  */
  assign level0_d1 = n1206; // (signal)
  /* fppowbf16.vhdl:2083:27  */
  assign level0_d2 = n1207; // (signal)
  /* fppowbf16.vhdl:2083:38  */
  assign level0_d3 = n1208; // (signal)
  /* fppowbf16.vhdl:2085:8  */
  assign level1 = n1183; // (signal)
  /* fppowbf16.vhdl:2085:16  */
  assign level1_d1 = n1209; // (signal)
  /* fppowbf16.vhdl:2087:8  */
  assign level2 = n1189; // (signal)
  /* fppowbf16.vhdl:2089:8  */
  assign level3 = n1195; // (signal)
  /* fppowbf16.vhdl:2091:8  */
  assign level4 = n1201; // (signal)
  /* fppowbf16.vhdl:2106:23  */
  assign n1181 = {level0_d3, 1'b0};
  /* fppowbf16.vhdl:2106:52  */
  assign n1182 = ps[0]; // extract
  /* fppowbf16.vhdl:2106:45  */
  assign n1183 = n1182 ? n1181 : n1185;
  /* fppowbf16.vhdl:2106:90  */
  assign n1185 = {1'b0, level0_d3};
  /* fppowbf16.vhdl:2107:23  */
  assign n1187 = {level1_d1, 2'b00};
  /* fppowbf16.vhdl:2107:55  */
  assign n1188 = ps_d1[1]; // extract
  /* fppowbf16.vhdl:2107:45  */
  assign n1189 = n1188 ? n1187 : n1191;
  /* fppowbf16.vhdl:2107:93  */
  assign n1191 = {2'b00, level1_d1};
  /* fppowbf16.vhdl:2108:20  */
  assign n1193 = {level2, 4'b0000};
  /* fppowbf16.vhdl:2108:52  */
  assign n1194 = ps_d1[2]; // extract
  /* fppowbf16.vhdl:2108:42  */
  assign n1195 = n1194 ? n1193 : n1197;
  /* fppowbf16.vhdl:2108:90  */
  assign n1197 = {4'b0000, level2};
  /* fppowbf16.vhdl:2109:20  */
  assign n1199 = {level3, 8'b00000000};
  /* fppowbf16.vhdl:2109:52  */
  assign n1200 = ps_d1[3]; // extract
  /* fppowbf16.vhdl:2109:42  */
  assign n1201 = n1200 ? n1199 : n1203;
  /* fppowbf16.vhdl:2109:90  */
  assign n1203 = {8'b00000000, level3};
  /* fppowbf16.vhdl:2110:15  */
  assign n1204 = level4[19:0]; // extract
  /* fppowbf16.vhdl:2096:10  */
  always @(posedge clk)
    n1205 <= ps;
  /* fppowbf16.vhdl:2096:10  */
  always @(posedge clk)
    n1206 <= level0;
  /* fppowbf16.vhdl:2096:10  */
  always @(posedge clk)
    n1207 <= level0_d1;
  /* fppowbf16.vhdl:2096:10  */
  always @(posedge clk)
    n1208 <= level0_d2;
  /* fppowbf16.vhdl:2096:10  */
  always @(posedge clk)
    n1209 <= level1;
endmodule

module lzoc_17_freq500_uid11
  (input  clk,
   input  [16:0] i,
   input  ozb,
   output [4:0] o);
  wire sozb;
  wire sozb_d1;
  wire sozb_d2;
  wire [30:0] level5;
  wire [30:0] level5_d1;
  wire digit4;
  wire digit4_d1;
  wire digit4_d2;
  wire [14:0] level4;
  wire [14:0] level4_d1;
  wire digit3;
  wire digit3_d1;
  wire [6:0] level3;
  wire digit2;
  wire [2:0] level2;
  wire [2:0] level2_d1;
  wire [2:0] z;
  wire [1:0] lowbits;
  wire [2:0] outhighbits;
  wire [2:0] outhighbits_d1;
  wire ozb_d1;
  wire ozb_d2;
  wire ozb_d3;
  wire n1083;
  wire n1084;
  wire n1085;
  wire n1086;
  wire n1087;
  wire n1088;
  wire n1089;
  wire n1090;
  wire n1091;
  wire n1092;
  wire n1093;
  wire n1094;
  wire n1095;
  wire n1096;
  wire [3:0] n1097;
  wire [3:0] n1098;
  wire [3:0] n1099;
  wire [1:0] n1100;
  wire [13:0] n1101;
  wire [30:0] n1102;
  wire [15:0] n1104;
  wire [3:0] n1105;
  wire [3:0] n1106;
  wire [3:0] n1107;
  wire [3:0] n1108;
  wire [15:0] n1109;
  wire n1110;
  wire n1111;
  wire [14:0] n1113;
  wire [14:0] n1114;
  wire [14:0] n1115;
  wire [7:0] n1117;
  wire [3:0] n1118;
  wire [3:0] n1119;
  wire [7:0] n1120;
  wire n1121;
  wire n1122;
  wire [6:0] n1124;
  wire [6:0] n1125;
  wire [6:0] n1126;
  wire [3:0] n1128;
  wire [3:0] n1129;
  wire n1130;
  wire n1131;
  wire [2:0] n1133;
  wire [2:0] n1134;
  wire [2:0] n1135;
  wire n1136;
  wire [2:0] n1137;
  wire [2:0] n1138;
  wire n1141;
  wire n1144;
  wire n1147;
  wire n1150;
  wire [3:0] n1152;
  reg [1:0] n1153;
  wire [1:0] n1154;
  wire [2:0] n1155;
  wire [4:0] n1157;
  reg n1158;
  reg n1159;
  reg [30:0] n1160;
  reg n1161;
  reg n1162;
  reg [14:0] n1163;
  reg n1164;
  reg [2:0] n1165;
  reg [2:0] n1166;
  reg n1167;
  reg n1168;
  reg n1169;
  assign o = n1157; //(module output)
  /* fppowbf16.vhdl:1986:8  */
  assign sozb = ozb; // (signal)
  /* fppowbf16.vhdl:1986:14  */
  assign sozb_d1 = n1158; // (signal)
  /* fppowbf16.vhdl:1986:23  */
  assign sozb_d2 = n1159; // (signal)
  /* fppowbf16.vhdl:1988:8  */
  assign level5 = n1102; // (signal)
  /* fppowbf16.vhdl:1988:16  */
  assign level5_d1 = n1160; // (signal)
  /* fppowbf16.vhdl:1990:8  */
  assign digit4 = n1111; // (signal)
  /* fppowbf16.vhdl:1990:16  */
  assign digit4_d1 = n1161; // (signal)
  /* fppowbf16.vhdl:1990:27  */
  assign digit4_d2 = n1162; // (signal)
  /* fppowbf16.vhdl:1992:8  */
  assign level4 = n1114; // (signal)
  /* fppowbf16.vhdl:1992:16  */
  assign level4_d1 = n1163; // (signal)
  /* fppowbf16.vhdl:1994:8  */
  assign digit3 = n1122; // (signal)
  /* fppowbf16.vhdl:1994:16  */
  assign digit3_d1 = n1164; // (signal)
  /* fppowbf16.vhdl:1996:8  */
  assign level3 = n1125; // (signal)
  /* fppowbf16.vhdl:1998:8  */
  assign digit2 = n1131; // (signal)
  /* fppowbf16.vhdl:2000:8  */
  assign level2 = n1134; // (signal)
  /* fppowbf16.vhdl:2000:16  */
  assign level2_d1 = n1165; // (signal)
  /* fppowbf16.vhdl:2002:8  */
  assign z = n1137; // (signal)
  /* fppowbf16.vhdl:2004:8  */
  assign lowbits = n1153; // (signal)
  /* fppowbf16.vhdl:2006:8  */
  assign outhighbits = n1155; // (signal)
  /* fppowbf16.vhdl:2006:21  */
  assign outhighbits_d1 = n1166; // (signal)
  /* fppowbf16.vhdl:2008:8  */
  assign ozb_d1 = n1167; // (signal)
  /* fppowbf16.vhdl:2008:16  */
  assign ozb_d2 = n1168; // (signal)
  /* fppowbf16.vhdl:2008:24  */
  assign ozb_d3 = n1169; // (signal)
  /* fppowbf16.vhdl:2030:34  */
  assign n1083 = ~sozb;
  /* fppowbf16.vhdl:2030:34  */
  assign n1084 = ~sozb;
  /* fppowbf16.vhdl:2030:34  */
  assign n1085 = ~sozb;
  /* fppowbf16.vhdl:2030:34  */
  assign n1086 = ~sozb;
  /* fppowbf16.vhdl:2030:34  */
  assign n1087 = ~sozb;
  /* fppowbf16.vhdl:2030:34  */
  assign n1088 = ~sozb;
  /* fppowbf16.vhdl:2030:34  */
  assign n1089 = ~sozb;
  /* fppowbf16.vhdl:2030:34  */
  assign n1090 = ~sozb;
  /* fppowbf16.vhdl:2030:34  */
  assign n1091 = ~sozb;
  /* fppowbf16.vhdl:2030:34  */
  assign n1092 = ~sozb;
  /* fppowbf16.vhdl:2030:34  */
  assign n1093 = ~sozb;
  /* fppowbf16.vhdl:2030:34  */
  assign n1094 = ~sozb;
  /* fppowbf16.vhdl:2030:34  */
  assign n1095 = ~sozb;
  /* fppowbf16.vhdl:2030:34  */
  assign n1096 = ~sozb;
  assign n1097 = {n1096, n1095, n1094, n1093};
  assign n1098 = {n1092, n1091, n1090, n1089};
  assign n1099 = {n1088, n1087, n1086, n1085};
  assign n1100 = {n1084, n1083};
  assign n1101 = {n1097, n1098, n1099, n1100};
  /* fppowbf16.vhdl:2030:16  */
  assign n1102 = {i, n1101};
  /* fppowbf16.vhdl:2032:28  */
  assign n1104 = level5[30:15]; // extract
  assign n1105 = {sozb, sozb, sozb, sozb};
  assign n1106 = {sozb, sozb, sozb, sozb};
  assign n1107 = {sozb, sozb, sozb, sozb};
  assign n1108 = {sozb, sozb, sozb, sozb};
  assign n1109 = {n1105, n1106, n1107, n1108};
  /* fppowbf16.vhdl:2032:43  */
  assign n1110 = n1104 == n1109;
  /* fppowbf16.vhdl:2032:17  */
  assign n1111 = n1110 ? 1'b1 : 1'b0;
  /* fppowbf16.vhdl:2033:22  */
  assign n1113 = level5_d1[14:0]; // extract
  /* fppowbf16.vhdl:2033:36  */
  assign n1114 = digit4_d1 ? n1113 : n1115;
  /* fppowbf16.vhdl:2033:69  */
  assign n1115 = level5_d1[30:16]; // extract
  /* fppowbf16.vhdl:2034:28  */
  assign n1117 = level4[14:7]; // extract
  assign n1118 = {sozb_d1, sozb_d1, sozb_d1, sozb_d1};
  assign n1119 = {sozb_d1, sozb_d1, sozb_d1, sozb_d1};
  assign n1120 = {n1118, n1119};
  /* fppowbf16.vhdl:2034:42  */
  assign n1121 = n1117 == n1120;
  /* fppowbf16.vhdl:2034:17  */
  assign n1122 = n1121 ? 1'b1 : 1'b0;
  /* fppowbf16.vhdl:2035:22  */
  assign n1124 = level4_d1[6:0]; // extract
  /* fppowbf16.vhdl:2035:35  */
  assign n1125 = digit3_d1 ? n1124 : n1126;
  /* fppowbf16.vhdl:2035:68  */
  assign n1126 = level4_d1[14:8]; // extract
  /* fppowbf16.vhdl:2036:28  */
  assign n1128 = level3[6:3]; // extract
  assign n1129 = {sozb_d2, sozb_d2, sozb_d2, sozb_d2};
  /* fppowbf16.vhdl:2036:41  */
  assign n1130 = n1128 == n1129;
  /* fppowbf16.vhdl:2036:17  */
  assign n1131 = n1130 ? 1'b1 : 1'b0;
  /* fppowbf16.vhdl:2037:19  */
  assign n1133 = level3[2:0]; // extract
  /* fppowbf16.vhdl:2037:32  */
  assign n1134 = digit2 ? n1133 : n1135;
  /* fppowbf16.vhdl:2037:59  */
  assign n1135 = level3[6:4]; // extract
  /* fppowbf16.vhdl:2039:30  */
  assign n1136 = ~ozb_d3;
  /* fppowbf16.vhdl:2039:19  */
  assign n1137 = n1136 ? level2_d1 : n1138;
  /* fppowbf16.vhdl:2039:41  */
  assign n1138 = ~level2_d1;
  /* fppowbf16.vhdl:2041:12  */
  assign n1141 = z == 3'b000;
  /* fppowbf16.vhdl:2042:12  */
  assign n1144 = z == 3'b001;
  /* fppowbf16.vhdl:2043:12  */
  assign n1147 = z == 3'b010;
  /* fppowbf16.vhdl:2044:12  */
  assign n1150 = z == 3'b011;
  assign n1152 = {n1150, n1147, n1144, n1141};
  /* fppowbf16.vhdl:2040:4  */
  always @*
    case (n1152)
      4'b1000: n1153 = 2'b01;
      4'b0100: n1153 = 2'b01;
      4'b0010: n1153 = 2'b10;
      4'b0001: n1153 = 2'b11;
      default: n1153 = 2'b00;
    endcase
  /* fppowbf16.vhdl:2046:29  */
  assign n1154 = {digit4_d2, digit3_d1};
  /* fppowbf16.vhdl:2046:50  */
  assign n1155 = {n1154, digit2};
  /* fppowbf16.vhdl:2047:24  */
  assign n1157 = {outhighbits_d1, lowbits};
  /* fppowbf16.vhdl:2013:10  */
  always @(posedge clk)
    n1158 <= sozb;
  /* fppowbf16.vhdl:2013:10  */
  always @(posedge clk)
    n1159 <= sozb_d1;
  /* fppowbf16.vhdl:2013:10  */
  always @(posedge clk)
    n1160 <= level5;
  /* fppowbf16.vhdl:2013:10  */
  always @(posedge clk)
    n1161 <= digit4;
  /* fppowbf16.vhdl:2013:10  */
  always @(posedge clk)
    n1162 <= digit4_d1;
  /* fppowbf16.vhdl:2013:10  */
  always @(posedge clk)
    n1163 <= level4;
  /* fppowbf16.vhdl:2013:10  */
  always @(posedge clk)
    n1164 <= digit3;
  /* fppowbf16.vhdl:2013:10  */
  always @(posedge clk)
    n1165 <= level2;
  /* fppowbf16.vhdl:2013:10  */
  always @(posedge clk)
    n1166 <= outhighbits;
  /* fppowbf16.vhdl:2013:10  */
  always @(posedge clk)
    n1167 <= ozb;
  /* fppowbf16.vhdl:2013:10  */
  always @(posedge clk)
    n1168 <= ozb_d1;
  /* fppowbf16.vhdl:2013:10  */
  always @(posedge clk)
    n1169 <= ozb_d2;
endmodule

module fpexp_8_7_freq500_uid71
  (input  clk,
   input  [28:0] x,
   output [17:0] r);
  wire [1:0] xexn;
  wire [1:0] xexn_d1;
  wire [1:0] xexn_d2;
  wire xsign;
  wire xsign_d1;
  wire xsign_d2;
  wire [7:0] xexpfield;
  wire [7:0] xexpfield_d1;
  wire [17:0] xfrac;
  wire [9:0] e0;
  wire [9:0] e0_d1;
  wire [9:0] e0_d2;
  wire [9:0] e0_d3;
  wire [9:0] e0_d4;
  wire [9:0] e0_d5;
  wire [9:0] e0_d6;
  wire [9:0] e0_d7;
  wire [9:0] e0_d8;
  wire [9:0] e0_d9;
  wire [9:0] e0_d10;
  wire [9:0] e0_d11;
  wire [9:0] e0_d12;
  wire [9:0] e0_d13;
  wire [9:0] e0_d14;
  wire [9:0] shiftval;
  wire resultwillbeone;
  wire resultwillbeone_d1;
  wire [18:0] mxu;
  wire [8:0] maxshift;
  wire [8:0] maxshift_d1;
  wire [8:0] maxshift_d2;
  wire [8:0] maxshift_d3;
  wire [8:0] maxshift_d4;
  wire [8:0] maxshift_d5;
  wire [8:0] maxshift_d6;
  wire [8:0] maxshift_d7;
  wire [8:0] maxshift_d8;
  wire [8:0] maxshift_d9;
  wire [8:0] maxshift_d10;
  wire [8:0] maxshift_d11;
  wire [8:0] maxshift_d12;
  wire [8:0] maxshift_d13;
  wire [8:0] maxshift_d14;
  wire overflow0;
  wire overflow0_d1;
  wire [4:0] shiftvalin;
  wire [34:0] fixx0;
  wire [16:0] ufixx;
  wire [12:0] expy;
  wire [8:0] k;
  wire neednonorm;
  wire [16:0] preroundbiassig;
  wire roundbit;
  wire [16:0] roundnormaddend;
  wire [16:0] roundedexpsigres;
  wire [16:0] roundedexpsig;
  wire ofl1;
  wire ofl2;
  wire ofl3;
  wire ofl;
  wire ufl1;
  wire ufl2;
  wire ufl3;
  wire ufl;
  wire [1:0] rexn;
  wire [1:0] n915;
  wire n916;
  wire [7:0] n917;
  wire [17:0] n918;
  wire [9:0] n921;
  wire [9:0] n922;
  wire n923;
  wire [18:0] n925;
  wire n927;
  wire n928;
  wire [8:0] n929;
  wire n930;
  wire n931;
  wire [4:0] n933;
  wire [34:0] mantissa_shift_n934;
  wire [16:0] n937;
  wire n938;
  wire [16:0] n939;
  wire [12:0] exp_helper_n941;
  wire [8:0] exp_helper_n942;
  wire n947;
  wire [6:0] n948;
  wire [16:0] n950;
  wire [16:0] n951;
  wire [6:0] n952;
  wire [16:0] n954;
  wire n955;
  wire n956;
  wire n957;
  wire n958;
  wire [9:0] n959;
  wire [15:0] n961;
  wire [16:0] n962;
  localparam n963 = 1'b0;
  wire [16:0] roundedexpsigoperandadder_n964;
  wire n968;
  wire [16:0] n969;
  wire n971;
  wire n972;
  wire n973;
  wire n974;
  wire n975;
  wire n976;
  wire n977;
  wire n978;
  wire n979;
  wire n980;
  wire n981;
  wire n982;
  wire n983;
  wire n984;
  wire n985;
  wire n986;
  wire n987;
  wire n988;
  wire n989;
  wire n990;
  wire n991;
  wire n992;
  wire n993;
  wire n994;
  wire n995;
  wire n996;
  wire n997;
  wire n998;
  wire n999;
  wire n1000;
  wire n1001;
  wire n1002;
  wire n1003;
  wire n1004;
  wire n1005;
  wire n1006;
  wire n1007;
  wire n1008;
  wire n1009;
  wire n1010;
  wire n1011;
  wire n1012;
  wire n1013;
  wire n1014;
  wire n1015;
  wire n1016;
  wire n1017;
  wire n1020;
  wire [1:0] n1021;
  wire [1:0] n1023;
  wire [1:0] n1025;
  wire [2:0] n1028;
  wire [14:0] n1029;
  wire [17:0] n1030;
  reg [1:0] n1031;
  reg [1:0] n1032;
  reg n1033;
  reg n1034;
  reg [7:0] n1035;
  reg [9:0] n1036;
  reg [9:0] n1037;
  reg [9:0] n1038;
  reg [9:0] n1039;
  reg [9:0] n1040;
  reg [9:0] n1041;
  reg [9:0] n1042;
  reg [9:0] n1043;
  reg [9:0] n1044;
  reg [9:0] n1045;
  reg [9:0] n1046;
  reg [9:0] n1047;
  reg [9:0] n1048;
  reg [9:0] n1049;
  reg n1050;
  reg [8:0] n1051;
  reg [8:0] n1052;
  reg [8:0] n1053;
  reg [8:0] n1054;
  reg [8:0] n1055;
  reg [8:0] n1056;
  reg [8:0] n1057;
  reg [8:0] n1058;
  reg [8:0] n1059;
  reg [8:0] n1060;
  reg [8:0] n1061;
  reg [8:0] n1062;
  reg [8:0] n1063;
  reg [8:0] n1064;
  reg n1065;
  assign r = n1030; //(module output)
  /* fppowbf16.vhdl:4807:8  */
  assign xexn = n915; // (signal)
  /* fppowbf16.vhdl:4807:14  */
  assign xexn_d1 = n1031; // (signal)
  /* fppowbf16.vhdl:4807:23  */
  assign xexn_d2 = n1032; // (signal)
  /* fppowbf16.vhdl:4809:8  */
  assign xsign = n916; // (signal)
  /* fppowbf16.vhdl:4809:15  */
  assign xsign_d1 = n1033; // (signal)
  /* fppowbf16.vhdl:4809:25  */
  assign xsign_d2 = n1034; // (signal)
  /* fppowbf16.vhdl:4811:8  */
  assign xexpfield = n917; // (signal)
  /* fppowbf16.vhdl:4811:19  */
  assign xexpfield_d1 = n1035; // (signal)
  /* fppowbf16.vhdl:4813:8  */
  assign xfrac = n918; // (signal)
  /* fppowbf16.vhdl:4815:8  */
  assign e0 = 10'b0001110101; // (signal)
  /* fppowbf16.vhdl:4815:12  */
  assign e0_d1 = n1036; // (signal)
  /* fppowbf16.vhdl:4815:19  */
  assign e0_d2 = n1037; // (signal)
  /* fppowbf16.vhdl:4815:26  */
  assign e0_d3 = n1038; // (signal)
  /* fppowbf16.vhdl:4815:33  */
  assign e0_d4 = n1039; // (signal)
  /* fppowbf16.vhdl:4815:40  */
  assign e0_d5 = n1040; // (signal)
  /* fppowbf16.vhdl:4815:47  */
  assign e0_d6 = n1041; // (signal)
  /* fppowbf16.vhdl:4815:54  */
  assign e0_d7 = n1042; // (signal)
  /* fppowbf16.vhdl:4815:61  */
  assign e0_d8 = n1043; // (signal)
  /* fppowbf16.vhdl:4815:68  */
  assign e0_d9 = n1044; // (signal)
  /* fppowbf16.vhdl:4815:75  */
  assign e0_d10 = n1045; // (signal)
  /* fppowbf16.vhdl:4815:83  */
  assign e0_d11 = n1046; // (signal)
  /* fppowbf16.vhdl:4815:91  */
  assign e0_d12 = n1047; // (signal)
  /* fppowbf16.vhdl:4815:99  */
  assign e0_d13 = n1048; // (signal)
  /* fppowbf16.vhdl:4815:107  */
  assign e0_d14 = n1049; // (signal)
  /* fppowbf16.vhdl:4817:8  */
  assign shiftval = n922; // (signal)
  /* fppowbf16.vhdl:4819:8  */
  assign resultwillbeone = n923; // (signal)
  /* fppowbf16.vhdl:4819:25  */
  assign resultwillbeone_d1 = n1050; // (signal)
  /* fppowbf16.vhdl:4821:8  */
  assign mxu = n925; // (signal)
  /* fppowbf16.vhdl:4823:8  */
  assign maxshift = 9'b000010000; // (signal)
  /* fppowbf16.vhdl:4823:18  */
  assign maxshift_d1 = n1051; // (signal)
  /* fppowbf16.vhdl:4823:31  */
  assign maxshift_d2 = n1052; // (signal)
  /* fppowbf16.vhdl:4823:44  */
  assign maxshift_d3 = n1053; // (signal)
  /* fppowbf16.vhdl:4823:57  */
  assign maxshift_d4 = n1054; // (signal)
  /* fppowbf16.vhdl:4823:70  */
  assign maxshift_d5 = n1055; // (signal)
  /* fppowbf16.vhdl:4823:83  */
  assign maxshift_d6 = n1056; // (signal)
  /* fppowbf16.vhdl:4823:96  */
  assign maxshift_d7 = n1057; // (signal)
  /* fppowbf16.vhdl:4823:109  */
  assign maxshift_d8 = n1058; // (signal)
  /* fppowbf16.vhdl:4823:122  */
  assign maxshift_d9 = n1059; // (signal)
  /* fppowbf16.vhdl:4823:135  */
  assign maxshift_d10 = n1060; // (signal)
  /* fppowbf16.vhdl:4823:149  */
  assign maxshift_d11 = n1061; // (signal)
  /* fppowbf16.vhdl:4823:163  */
  assign maxshift_d12 = n1062; // (signal)
  /* fppowbf16.vhdl:4823:177  */
  assign maxshift_d13 = n1063; // (signal)
  /* fppowbf16.vhdl:4823:191  */
  assign maxshift_d14 = n1064; // (signal)
  /* fppowbf16.vhdl:4825:8  */
  assign overflow0 = n931; // (signal)
  /* fppowbf16.vhdl:4825:19  */
  assign overflow0_d1 = n1065; // (signal)
  /* fppowbf16.vhdl:4827:8  */
  assign shiftvalin = n933; // (signal)
  /* fppowbf16.vhdl:4829:8  */
  assign fixx0 = mantissa_shift_n934; // (signal)
  /* fppowbf16.vhdl:4831:8  */
  assign ufixx = n939; // (signal)
  /* fppowbf16.vhdl:4833:8  */
  assign expy = exp_helper_n941; // (signal)
  /* fppowbf16.vhdl:4835:8  */
  assign k = exp_helper_n942; // (signal)
  /* fppowbf16.vhdl:4837:8  */
  assign neednonorm = n947; // (signal)
  /* fppowbf16.vhdl:4839:8  */
  assign preroundbiassig = n951; // (signal)
  /* fppowbf16.vhdl:4841:8  */
  assign roundbit = n956; // (signal)
  /* fppowbf16.vhdl:4843:8  */
  assign roundnormaddend = n962; // (signal)
  /* fppowbf16.vhdl:4845:8  */
  assign roundedexpsigres = roundedexpsigoperandadder_n964; // (signal)
  /* fppowbf16.vhdl:4847:8  */
  assign roundedexpsig = n969; // (signal)
  /* fppowbf16.vhdl:4849:8  */
  assign ofl1 = n977; // (signal)
  /* fppowbf16.vhdl:4851:8  */
  assign ofl2 = n988; // (signal)
  /* fppowbf16.vhdl:4853:8  */
  assign ofl3 = n994; // (signal)
  /* fppowbf16.vhdl:4855:8  */
  assign ofl = n996; // (signal)
  /* fppowbf16.vhdl:4857:8  */
  assign ufl1 = n1004; // (signal)
  /* fppowbf16.vhdl:4859:8  */
  assign ufl2 = n1009; // (signal)
  /* fppowbf16.vhdl:4861:8  */
  assign ufl3 = n1015; // (signal)
  /* fppowbf16.vhdl:4863:8  */
  assign ufl = n1017; // (signal)
  /* fppowbf16.vhdl:4865:8  */
  assign rexn = n1021; // (signal)
  /* fppowbf16.vhdl:4912:13  */
  assign n915 = x[28:27]; // extract
  /* fppowbf16.vhdl:4913:14  */
  assign n916 = x[26]; // extract
  /* fppowbf16.vhdl:4914:18  */
  assign n917 = x[25:18]; // extract
  /* fppowbf16.vhdl:4915:23  */
  assign n918 = x[17:0]; // extract
  /* fppowbf16.vhdl:4917:22  */
  assign n921 = {2'b00, xexpfield_d1};
  /* fppowbf16.vhdl:4917:38  */
  assign n922 = n921 - e0_d14;
  /* fppowbf16.vhdl:4919:31  */
  assign n923 = shiftval[9]; // extract
  /* fppowbf16.vhdl:4921:15  */
  assign n925 = {1'b1, xfrac};
  /* fppowbf16.vhdl:4924:29  */
  assign n927 = shiftval[9]; // extract
  /* fppowbf16.vhdl:4924:17  */
  assign n928 = ~n927;
  /* fppowbf16.vhdl:4924:49  */
  assign n929 = shiftval[8:0]; // extract
  /* fppowbf16.vhdl:4924:63  */
  assign n930 = $unsigned(n929) > $unsigned(maxshift_d14);
  /* fppowbf16.vhdl:4924:36  */
  assign n931 = n930 ? n928 : 1'b0;
  /* fppowbf16.vhdl:4925:26  */
  assign n933 = shiftval[4:0]; // extract
  /* fppowbf16.vhdl:4926:4  */
  leftshifter19_by_max_16_freq500_uid73 mantissa_shift (
    .clk(clk),
    .x(mxu),
    .s(shiftvalin),
    .r(mantissa_shift_n934));
  /* fppowbf16.vhdl:4931:28  */
  assign n937 = fixx0[34:18]; // extract
  /* fppowbf16.vhdl:4931:67  */
  assign n938 = ~resultwillbeone_d1;
  /* fppowbf16.vhdl:4931:44  */
  assign n939 = n938 ? n937 : 17'b00000000000000000;
  /* fppowbf16.vhdl:4932:4  */
  exp_8_7_freq500_uid75 exp_helper (
    .clk(clk),
    .ufixx_i(ufixx),
    .xsign(xsign),
    .expy(exp_helper_n941),
    .k(exp_helper_n942));
  /* fppowbf16.vhdl:4938:22  */
  assign n947 = expy[12]; // extract
  /* fppowbf16.vhdl:4940:63  */
  assign n948 = expy[11:5]; // extract
  /* fppowbf16.vhdl:4940:57  */
  assign n950 = {10'b0001111111, n948};
  /* fppowbf16.vhdl:4940:77  */
  assign n951 = neednonorm ? n950 : n954;
  /* fppowbf16.vhdl:4941:52  */
  assign n952 = expy[10:4]; // extract
  /* fppowbf16.vhdl:4941:46  */
  assign n954 = {10'b0001111110, n952};
  /* fppowbf16.vhdl:4942:20  */
  assign n955 = expy[4]; // extract
  /* fppowbf16.vhdl:4942:25  */
  assign n956 = neednonorm ? n955 : n957;
  /* fppowbf16.vhdl:4942:59  */
  assign n957 = expy[3]; // extract
  /* fppowbf16.vhdl:4943:24  */
  assign n958 = k[8]; // extract
  /* fppowbf16.vhdl:4943:28  */
  assign n959 = {n958, k};
  /* fppowbf16.vhdl:4943:32  */
  assign n961 = {n959, 6'b000000};
  /* fppowbf16.vhdl:4943:54  */
  assign n962 = {n961, roundbit};
  /* fppowbf16.vhdl:4944:4  */
  intadder_17_freq500_uid107 roundedexpsigoperandadder (
    .clk(clk),
    .x(preroundbiassig),
    .y(roundnormaddend),
    .cin(n963),
    .r(roundedexpsigoperandadder_n964));
  /* fppowbf16.vhdl:4950:47  */
  assign n968 = xexn == 2'b01;
  /* fppowbf16.vhdl:4950:38  */
  assign n969 = n968 ? roundedexpsigres : 17'b00011111110000000;
  /* fppowbf16.vhdl:4951:12  */
  assign n971 = ~xsign_d2;
  /* fppowbf16.vhdl:4951:25  */
  assign n972 = n971 & overflow0_d1;
  /* fppowbf16.vhdl:4951:58  */
  assign n973 = xexn_d2[1]; // extract
  /* fppowbf16.vhdl:4951:47  */
  assign n974 = ~n973;
  /* fppowbf16.vhdl:4951:73  */
  assign n975 = xexn_d2[0]; // extract
  /* fppowbf16.vhdl:4951:62  */
  assign n976 = n974 & n975;
  /* fppowbf16.vhdl:4951:42  */
  assign n977 = n972 & n976;
  /* fppowbf16.vhdl:4952:12  */
  assign n978 = ~xsign;
  /* fppowbf16.vhdl:4952:40  */
  assign n979 = roundedexpsig[15]; // extract
  /* fppowbf16.vhdl:4952:69  */
  assign n980 = roundedexpsig[16]; // extract
  /* fppowbf16.vhdl:4952:52  */
  assign n981 = ~n980;
  /* fppowbf16.vhdl:4952:48  */
  assign n982 = n979 & n981;
  /* fppowbf16.vhdl:4952:22  */
  assign n983 = n978 & n982;
  /* fppowbf16.vhdl:4952:93  */
  assign n984 = xexn[1]; // extract
  /* fppowbf16.vhdl:4952:85  */
  assign n985 = ~n984;
  /* fppowbf16.vhdl:4952:105  */
  assign n986 = xexn[0]; // extract
  /* fppowbf16.vhdl:4952:97  */
  assign n987 = n985 & n986;
  /* fppowbf16.vhdl:4952:80  */
  assign n988 = n983 & n987;
  /* fppowbf16.vhdl:4953:12  */
  assign n989 = ~xsign;
  /* fppowbf16.vhdl:4953:30  */
  assign n990 = xexn[1]; // extract
  /* fppowbf16.vhdl:4953:22  */
  assign n991 = n989 & n990;
  /* fppowbf16.vhdl:4953:46  */
  assign n992 = xexn[0]; // extract
  /* fppowbf16.vhdl:4953:38  */
  assign n993 = ~n992;
  /* fppowbf16.vhdl:4953:34  */
  assign n994 = n991 & n993;
  /* fppowbf16.vhdl:4954:16  */
  assign n995 = ofl1 | ofl2;
  /* fppowbf16.vhdl:4954:24  */
  assign n996 = n995 | ofl3;
  /* fppowbf16.vhdl:4955:26  */
  assign n997 = roundedexpsig[15]; // extract
  /* fppowbf16.vhdl:4955:51  */
  assign n998 = roundedexpsig[16]; // extract
  /* fppowbf16.vhdl:4955:34  */
  assign n999 = n997 & n998;
  /* fppowbf16.vhdl:4955:76  */
  assign n1000 = xexn[1]; // extract
  /* fppowbf16.vhdl:4955:68  */
  assign n1001 = ~n1000;
  /* fppowbf16.vhdl:4955:88  */
  assign n1002 = xexn[0]; // extract
  /* fppowbf16.vhdl:4955:80  */
  assign n1003 = n1001 & n1002;
  /* fppowbf16.vhdl:4955:63  */
  assign n1004 = n999 & n1003;
  /* fppowbf16.vhdl:4956:26  */
  assign n1005 = xexn[1]; // extract
  /* fppowbf16.vhdl:4956:18  */
  assign n1006 = xsign & n1005;
  /* fppowbf16.vhdl:4956:42  */
  assign n1007 = xexn[0]; // extract
  /* fppowbf16.vhdl:4956:34  */
  assign n1008 = ~n1007;
  /* fppowbf16.vhdl:4956:30  */
  assign n1009 = n1006 & n1008;
  /* fppowbf16.vhdl:4957:21  */
  assign n1010 = xsign_d1 & overflow0;
  /* fppowbf16.vhdl:4957:52  */
  assign n1011 = xexn_d1[1]; // extract
  /* fppowbf16.vhdl:4957:41  */
  assign n1012 = ~n1011;
  /* fppowbf16.vhdl:4957:67  */
  assign n1013 = xexn_d1[0]; // extract
  /* fppowbf16.vhdl:4957:56  */
  assign n1014 = n1012 & n1013;
  /* fppowbf16.vhdl:4957:36  */
  assign n1015 = n1010 & n1014;
  /* fppowbf16.vhdl:4958:16  */
  assign n1016 = ufl1 | ufl2;
  /* fppowbf16.vhdl:4958:24  */
  assign n1017 = n1016 | ufl3;
  /* fppowbf16.vhdl:4959:27  */
  assign n1020 = xexn == 2'b11;
  /* fppowbf16.vhdl:4959:17  */
  assign n1021 = n1020 ? 2'b11 : n1023;
  /* fppowbf16.vhdl:4960:7  */
  assign n1023 = ofl ? 2'b10 : n1025;
  /* fppowbf16.vhdl:4961:7  */
  assign n1025 = ufl ? 2'b00 : 2'b01;
  /* fppowbf16.vhdl:4963:14  */
  assign n1028 = {rexn, 1'b0};
  /* fppowbf16.vhdl:4963:35  */
  assign n1029 = roundedexpsig[14:0]; // extract
  /* fppowbf16.vhdl:4963:20  */
  assign n1030 = {n1028, n1029};
  /* fppowbf16.vhdl:4874:10  */
  always @(posedge clk)
    n1031 <= xexn;
  /* fppowbf16.vhdl:4874:10  */
  always @(posedge clk)
    n1032 <= xexn_d1;
  /* fppowbf16.vhdl:4874:10  */
  always @(posedge clk)
    n1033 <= xsign;
  /* fppowbf16.vhdl:4874:10  */
  always @(posedge clk)
    n1034 <= xsign_d1;
  /* fppowbf16.vhdl:4874:10  */
  always @(posedge clk)
    n1035 <= xexpfield;
  /* fppowbf16.vhdl:4874:10  */
  always @(posedge clk)
    n1036 <= e0;
  /* fppowbf16.vhdl:4874:10  */
  always @(posedge clk)
    n1037 <= e0_d1;
  /* fppowbf16.vhdl:4874:10  */
  always @(posedge clk)
    n1038 <= e0_d2;
  /* fppowbf16.vhdl:4874:10  */
  always @(posedge clk)
    n1039 <= e0_d3;
  /* fppowbf16.vhdl:4874:10  */
  always @(posedge clk)
    n1040 <= e0_d4;
  /* fppowbf16.vhdl:4874:10  */
  always @(posedge clk)
    n1041 <= e0_d5;
  /* fppowbf16.vhdl:4874:10  */
  always @(posedge clk)
    n1042 <= e0_d6;
  /* fppowbf16.vhdl:4874:10  */
  always @(posedge clk)
    n1043 <= e0_d7;
  /* fppowbf16.vhdl:4874:10  */
  always @(posedge clk)
    n1044 <= e0_d8;
  /* fppowbf16.vhdl:4874:10  */
  always @(posedge clk)
    n1045 <= e0_d9;
  /* fppowbf16.vhdl:4874:10  */
  always @(posedge clk)
    n1046 <= e0_d10;
  /* fppowbf16.vhdl:4874:10  */
  always @(posedge clk)
    n1047 <= e0_d11;
  /* fppowbf16.vhdl:4874:10  */
  always @(posedge clk)
    n1048 <= e0_d12;
  /* fppowbf16.vhdl:4874:10  */
  always @(posedge clk)
    n1049 <= e0_d13;
  /* fppowbf16.vhdl:4874:10  */
  always @(posedge clk)
    n1050 <= resultwillbeone;
  /* fppowbf16.vhdl:4874:10  */
  always @(posedge clk)
    n1051 <= maxshift;
  /* fppowbf16.vhdl:4874:10  */
  always @(posedge clk)
    n1052 <= maxshift_d1;
  /* fppowbf16.vhdl:4874:10  */
  always @(posedge clk)
    n1053 <= maxshift_d2;
  /* fppowbf16.vhdl:4874:10  */
  always @(posedge clk)
    n1054 <= maxshift_d3;
  /* fppowbf16.vhdl:4874:10  */
  always @(posedge clk)
    n1055 <= maxshift_d4;
  /* fppowbf16.vhdl:4874:10  */
  always @(posedge clk)
    n1056 <= maxshift_d5;
  /* fppowbf16.vhdl:4874:10  */
  always @(posedge clk)
    n1057 <= maxshift_d6;
  /* fppowbf16.vhdl:4874:10  */
  always @(posedge clk)
    n1058 <= maxshift_d7;
  /* fppowbf16.vhdl:4874:10  */
  always @(posedge clk)
    n1059 <= maxshift_d8;
  /* fppowbf16.vhdl:4874:10  */
  always @(posedge clk)
    n1060 <= maxshift_d9;
  /* fppowbf16.vhdl:4874:10  */
  always @(posedge clk)
    n1061 <= maxshift_d10;
  /* fppowbf16.vhdl:4874:10  */
  always @(posedge clk)
    n1062 <= maxshift_d11;
  /* fppowbf16.vhdl:4874:10  */
  always @(posedge clk)
    n1063 <= maxshift_d12;
  /* fppowbf16.vhdl:4874:10  */
  always @(posedge clk)
    n1064 <= maxshift_d13;
  /* fppowbf16.vhdl:4874:10  */
  always @(posedge clk)
    n1065 <= overflow0;
endmodule

module fpmult_8_17_uid62_freq500_uid63
  (input  clk,
   input  [27:0] x,
   input  [17:0] y,
   output [28:0] r);
  wire sign;
  wire sign_d1;
  wire sign_d2;
  wire [7:0] expx;
  wire [7:0] expx_d1;
  wire [7:0] expy;
  wire [7:0] expy_d1;
  wire [7:0] expy_d2;
  wire [7:0] expy_d3;
  wire [7:0] expy_d4;
  wire [7:0] expy_d5;
  wire [7:0] expy_d6;
  wire [7:0] expy_d7;
  wire [7:0] expy_d8;
  wire [7:0] expy_d9;
  wire [7:0] expy_d10;
  wire [7:0] expy_d11;
  wire [7:0] expy_d12;
  wire [9:0] expsumpresub;
  wire [9:0] expsumpresub_d1;
  wire [9:0] bias;
  wire [9:0] bias_d1;
  wire [9:0] bias_d2;
  wire [9:0] bias_d3;
  wire [9:0] bias_d4;
  wire [9:0] bias_d5;
  wire [9:0] bias_d6;
  wire [9:0] bias_d7;
  wire [9:0] bias_d8;
  wire [9:0] bias_d9;
  wire [9:0] bias_d10;
  wire [9:0] bias_d11;
  wire [9:0] bias_d12;
  wire [9:0] bias_d13;
  wire [9:0] expsum;
  wire [17:0] sigx;
  wire [7:0] sigy;
  wire [20:0] sigprod;
  wire [20:0] sigprod_d1;
  wire [3:0] excsel;
  wire [1:0] exc;
  wire [1:0] exc_d1;
  wire [1:0] exc_d2;
  wire norm;
  wire norm_d1;
  wire norm_d2;
  wire [9:0] exppostnorm;
  wire [20:0] sigprodext;
  wire [20:0] sigprodext_d1;
  wire [27:0] expsig;
  wire round;
  wire [27:0] expsigpostround;
  wire [1:0] excpostnorm;
  wire [1:0] finalexc;
  wire [17:0] y_d1;
  wire [17:0] y_d2;
  wire [17:0] y_d3;
  wire [17:0] y_d4;
  wire [17:0] y_d5;
  wire [17:0] y_d6;
  wire [17:0] y_d7;
  wire [17:0] y_d8;
  wire [17:0] y_d9;
  wire [17:0] y_d10;
  wire [17:0] y_d11;
  wire n735;
  wire n736;
  wire n737;
  wire [7:0] n738;
  wire [7:0] n739;
  wire [9:0] n741;
  wire [9:0] n743;
  wire [9:0] n744;
  wire [9:0] n746;
  wire [16:0] n747;
  wire [17:0] n749;
  wire [6:0] n750;
  wire [7:0] n752;
  wire [20:0] significandmultiplication_n753;
  wire [1:0] n756;
  wire [1:0] n757;
  wire [3:0] n758;
  wire n761;
  wire n763;
  wire n764;
  wire n766;
  wire n767;
  wire n770;
  wire n773;
  wire n775;
  wire n776;
  wire n778;
  wire n779;
  wire [2:0] n781;
  reg [1:0] n782;
  wire n783;
  wire [9:0] n785;
  wire [9:0] n786;
  wire [19:0] n787;
  wire [20:0] n789;
  wire [20:0] n790;
  wire [18:0] n791;
  wire [20:0] n793;
  wire [17:0] n794;
  wire [27:0] n795;
  localparam [27:0] n797 = 28'b0000000000000000000000000000;
  wire [27:0] roundingadder_n798;
  wire [1:0] n801;
  wire n804;
  wire n807;
  wire n810;
  wire n812;
  wire n813;
  wire [2:0] n815;
  reg [1:0] n816;
  wire n818;
  wire n820;
  wire n821;
  wire n823;
  wire n824;
  reg [1:0] n825;
  wire [2:0] n826;
  wire [25:0] n827;
  wire [28:0] n828;
  reg n829;
  reg n830;
  reg [7:0] n831;
  reg [7:0] n832;
  reg [7:0] n833;
  reg [7:0] n834;
  reg [7:0] n835;
  reg [7:0] n836;
  reg [7:0] n837;
  reg [7:0] n838;
  reg [7:0] n839;
  reg [7:0] n840;
  reg [7:0] n841;
  reg [7:0] n842;
  reg [7:0] n843;
  reg [9:0] n844;
  reg [9:0] n845;
  reg [9:0] n846;
  reg [9:0] n847;
  reg [9:0] n848;
  reg [9:0] n849;
  reg [9:0] n850;
  reg [9:0] n851;
  reg [9:0] n852;
  reg [9:0] n853;
  reg [9:0] n854;
  reg [9:0] n855;
  reg [9:0] n856;
  reg [9:0] n857;
  reg [20:0] n858;
  reg [1:0] n859;
  reg [1:0] n860;
  reg n861;
  reg n862;
  reg [20:0] n863;
  reg [17:0] n864;
  reg [17:0] n865;
  reg [17:0] n866;
  reg [17:0] n867;
  reg [17:0] n868;
  reg [17:0] n869;
  reg [17:0] n870;
  reg [17:0] n871;
  reg [17:0] n872;
  reg [17:0] n873;
  reg [17:0] n874;
  assign r = n828; //(module output)
  /* fppowbf16.vhdl:3838:8  */
  assign sign = n737; // (signal)
  /* fppowbf16.vhdl:3838:14  */
  assign sign_d1 = n829; // (signal)
  /* fppowbf16.vhdl:3838:23  */
  assign sign_d2 = n830; // (signal)
  /* fppowbf16.vhdl:3840:8  */
  assign expx = n738; // (signal)
  /* fppowbf16.vhdl:3840:14  */
  assign expx_d1 = n831; // (signal)
  /* fppowbf16.vhdl:3842:8  */
  assign expy = n739; // (signal)
  /* fppowbf16.vhdl:3842:14  */
  assign expy_d1 = n832; // (signal)
  /* fppowbf16.vhdl:3842:23  */
  assign expy_d2 = n833; // (signal)
  /* fppowbf16.vhdl:3842:32  */
  assign expy_d3 = n834; // (signal)
  /* fppowbf16.vhdl:3842:41  */
  assign expy_d4 = n835; // (signal)
  /* fppowbf16.vhdl:3842:50  */
  assign expy_d5 = n836; // (signal)
  /* fppowbf16.vhdl:3842:59  */
  assign expy_d6 = n837; // (signal)
  /* fppowbf16.vhdl:3842:68  */
  assign expy_d7 = n838; // (signal)
  /* fppowbf16.vhdl:3842:77  */
  assign expy_d8 = n839; // (signal)
  /* fppowbf16.vhdl:3842:86  */
  assign expy_d9 = n840; // (signal)
  /* fppowbf16.vhdl:3842:95  */
  assign expy_d10 = n841; // (signal)
  /* fppowbf16.vhdl:3842:105  */
  assign expy_d11 = n842; // (signal)
  /* fppowbf16.vhdl:3842:115  */
  assign expy_d12 = n843; // (signal)
  /* fppowbf16.vhdl:3844:8  */
  assign expsumpresub = n744; // (signal)
  /* fppowbf16.vhdl:3844:22  */
  assign expsumpresub_d1 = n844; // (signal)
  /* fppowbf16.vhdl:3846:8  */
  assign bias = 10'b0001111111; // (signal)
  /* fppowbf16.vhdl:3846:14  */
  assign bias_d1 = n845; // (signal)
  /* fppowbf16.vhdl:3846:23  */
  assign bias_d2 = n846; // (signal)
  /* fppowbf16.vhdl:3846:32  */
  assign bias_d3 = n847; // (signal)
  /* fppowbf16.vhdl:3846:41  */
  assign bias_d4 = n848; // (signal)
  /* fppowbf16.vhdl:3846:50  */
  assign bias_d5 = n849; // (signal)
  /* fppowbf16.vhdl:3846:59  */
  assign bias_d6 = n850; // (signal)
  /* fppowbf16.vhdl:3846:68  */
  assign bias_d7 = n851; // (signal)
  /* fppowbf16.vhdl:3846:77  */
  assign bias_d8 = n852; // (signal)
  /* fppowbf16.vhdl:3846:86  */
  assign bias_d9 = n853; // (signal)
  /* fppowbf16.vhdl:3846:95  */
  assign bias_d10 = n854; // (signal)
  /* fppowbf16.vhdl:3846:105  */
  assign bias_d11 = n855; // (signal)
  /* fppowbf16.vhdl:3846:115  */
  assign bias_d12 = n856; // (signal)
  /* fppowbf16.vhdl:3846:125  */
  assign bias_d13 = n857; // (signal)
  /* fppowbf16.vhdl:3848:8  */
  assign expsum = n746; // (signal)
  /* fppowbf16.vhdl:3850:8  */
  assign sigx = n749; // (signal)
  /* fppowbf16.vhdl:3852:8  */
  assign sigy = n752; // (signal)
  /* fppowbf16.vhdl:3854:8  */
  assign sigprod = significandmultiplication_n753; // (signal)
  /* fppowbf16.vhdl:3854:17  */
  assign sigprod_d1 = n858; // (signal)
  /* fppowbf16.vhdl:3856:8  */
  assign excsel = n758; // (signal)
  /* fppowbf16.vhdl:3858:8  */
  assign exc = n782; // (signal)
  /* fppowbf16.vhdl:3858:13  */
  assign exc_d1 = n859; // (signal)
  /* fppowbf16.vhdl:3858:21  */
  assign exc_d2 = n860; // (signal)
  /* fppowbf16.vhdl:3860:8  */
  assign norm = n783; // (signal)
  /* fppowbf16.vhdl:3860:14  */
  assign norm_d1 = n861; // (signal)
  /* fppowbf16.vhdl:3860:23  */
  assign norm_d2 = n862; // (signal)
  /* fppowbf16.vhdl:3862:8  */
  assign exppostnorm = n786; // (signal)
  /* fppowbf16.vhdl:3864:8  */
  assign sigprodext = n790; // (signal)
  /* fppowbf16.vhdl:3864:20  */
  assign sigprodext_d1 = n863; // (signal)
  /* fppowbf16.vhdl:3866:8  */
  assign expsig = n795; // (signal)
  /* fppowbf16.vhdl:3868:8  */
  assign round = 1'b1; // (signal)
  /* fppowbf16.vhdl:3870:8  */
  assign expsigpostround = roundingadder_n798; // (signal)
  /* fppowbf16.vhdl:3872:8  */
  assign excpostnorm = n816; // (signal)
  /* fppowbf16.vhdl:3874:8  */
  assign finalexc = n825; // (signal)
  /* fppowbf16.vhdl:3876:8  */
  assign y_d1 = n864; // (signal)
  /* fppowbf16.vhdl:3876:14  */
  assign y_d2 = n865; // (signal)
  /* fppowbf16.vhdl:3876:20  */
  assign y_d3 = n866; // (signal)
  /* fppowbf16.vhdl:3876:26  */
  assign y_d4 = n867; // (signal)
  /* fppowbf16.vhdl:3876:32  */
  assign y_d5 = n868; // (signal)
  /* fppowbf16.vhdl:3876:38  */
  assign y_d6 = n869; // (signal)
  /* fppowbf16.vhdl:3876:44  */
  assign y_d7 = n870; // (signal)
  /* fppowbf16.vhdl:3876:50  */
  assign y_d8 = n871; // (signal)
  /* fppowbf16.vhdl:3876:56  */
  assign y_d9 = n872; // (signal)
  /* fppowbf16.vhdl:3876:62  */
  assign y_d10 = n873; // (signal)
  /* fppowbf16.vhdl:3876:69  */
  assign y_d11 = n874; // (signal)
  /* fppowbf16.vhdl:3930:13  */
  assign n735 = x[25]; // extract
  /* fppowbf16.vhdl:3930:27  */
  assign n736 = y_d11[15]; // extract
  /* fppowbf16.vhdl:3930:18  */
  assign n737 = n735 ^ n736;
  /* fppowbf16.vhdl:3931:13  */
  assign n738 = x[24:17]; // extract
  /* fppowbf16.vhdl:3932:13  */
  assign n739 = y[14:7]; // extract
  /* fppowbf16.vhdl:3933:26  */
  assign n741 = {2'b00, expx_d1};
  /* fppowbf16.vhdl:3933:45  */
  assign n743 = {2'b00, expy_d12};
  /* fppowbf16.vhdl:3933:37  */
  assign n744 = n741 + n743;
  /* fppowbf16.vhdl:3935:30  */
  assign n746 = expsumpresub_d1 - bias_d13;
  /* fppowbf16.vhdl:3936:19  */
  assign n747 = x[16:0]; // extract
  /* fppowbf16.vhdl:3936:16  */
  assign n749 = {1'b1, n747};
  /* fppowbf16.vhdl:3937:19  */
  assign n750 = y[6:0]; // extract
  /* fppowbf16.vhdl:3937:16  */
  assign n752 = {1'b1, n750};
  /* fppowbf16.vhdl:3938:4  */
  intmultiplier_18x8_21_freq500_uid65 significandmultiplication (
    .clk(clk),
    .x(sigx),
    .y(sigy),
    .r(significandmultiplication_n753));
  /* fppowbf16.vhdl:3943:15  */
  assign n756 = x[27:26]; // extract
  /* fppowbf16.vhdl:3943:37  */
  assign n757 = y_d11[17:16]; // extract
  /* fppowbf16.vhdl:3943:30  */
  assign n758 = {n756, n757};
  /* fppowbf16.vhdl:3945:16  */
  assign n761 = excsel == 4'b0000;
  /* fppowbf16.vhdl:3945:29  */
  assign n763 = excsel == 4'b0001;
  /* fppowbf16.vhdl:3945:29  */
  assign n764 = n761 | n763;
  /* fppowbf16.vhdl:3945:38  */
  assign n766 = excsel == 4'b0100;
  /* fppowbf16.vhdl:3945:38  */
  assign n767 = n764 | n766;
  /* fppowbf16.vhdl:3946:16  */
  assign n770 = excsel == 4'b0101;
  /* fppowbf16.vhdl:3947:16  */
  assign n773 = excsel == 4'b0110;
  /* fppowbf16.vhdl:3947:28  */
  assign n775 = excsel == 4'b1001;
  /* fppowbf16.vhdl:3947:28  */
  assign n776 = n773 | n775;
  /* fppowbf16.vhdl:3947:37  */
  assign n778 = excsel == 4'b1010;
  /* fppowbf16.vhdl:3947:37  */
  assign n779 = n776 | n778;
  assign n781 = {n779, n770, n767};
  /* fppowbf16.vhdl:3944:4  */
  always @*
    case (n781)
      3'b100: n782 = 2'b10;
      3'b010: n782 = 2'b01;
      3'b001: n782 = 2'b00;
      default: n782 = 2'b11;
    endcase
  /* fppowbf16.vhdl:3949:19  */
  assign n783 = sigprod[20]; // extract
  /* fppowbf16.vhdl:3951:41  */
  assign n785 = {9'b000000000, norm_d2};
  /* fppowbf16.vhdl:3951:26  */
  assign n786 = expsum + n785;
  /* fppowbf16.vhdl:3953:28  */
  assign n787 = sigprod_d1[19:0]; // extract
  /* fppowbf16.vhdl:3953:42  */
  assign n789 = {n787, 1'b0};
  /* fppowbf16.vhdl:3953:48  */
  assign n790 = norm_d1 ? n789 : n793;
  /* fppowbf16.vhdl:3954:36  */
  assign n791 = sigprod_d1[18:0]; // extract
  /* fppowbf16.vhdl:3954:50  */
  assign n793 = {n791, 2'b00};
  /* fppowbf16.vhdl:3955:41  */
  assign n794 = sigprodext_d1[20:3]; // extract
  /* fppowbf16.vhdl:3955:26  */
  assign n795 = {exppostnorm, n794};
  /* fppowbf16.vhdl:3957:4  */
  intadder_28_freq500_uid69 roundingadder (
    .clk(clk),
    .x(expsig),
    .y(n797),
    .cin(round),
    .r(roundingadder_n798));
  /* fppowbf16.vhdl:3963:24  */
  assign n801 = expsigpostround[27:26]; // extract
  /* fppowbf16.vhdl:3964:26  */
  assign n804 = n801 == 2'b00;
  /* fppowbf16.vhdl:3965:49  */
  assign n807 = n801 == 2'b01;
  /* fppowbf16.vhdl:3966:49  */
  assign n810 = n801 == 2'b11;
  /* fppowbf16.vhdl:3966:58  */
  assign n812 = n801 == 2'b10;
  /* fppowbf16.vhdl:3966:58  */
  assign n813 = n810 | n812;
  assign n815 = {n813, n807, n804};
  /* fppowbf16.vhdl:3963:4  */
  always @*
    case (n815)
      3'b100: n816 = 2'b00;
      3'b010: n816 = 2'b10;
      3'b001: n816 = 2'b01;
      default: n816 = 2'b11;
    endcase
  /* fppowbf16.vhdl:3969:23  */
  assign n818 = exc_d2 == 2'b11;
  /* fppowbf16.vhdl:3969:33  */
  assign n820 = exc_d2 == 2'b10;
  /* fppowbf16.vhdl:3969:33  */
  assign n821 = n818 | n820;
  /* fppowbf16.vhdl:3969:38  */
  assign n823 = exc_d2 == 2'b00;
  /* fppowbf16.vhdl:3969:38  */
  assign n824 = n821 | n823;
  /* fppowbf16.vhdl:3968:4  */
  always @*
    case (n824)
      1'b1: n825 = exc_d2;
      default: n825 = excpostnorm;
    endcase
  /* fppowbf16.vhdl:3971:18  */
  assign n826 = {finalexc, sign_d2};
  /* fppowbf16.vhdl:3971:45  */
  assign n827 = expsigpostround[25:0]; // extract
  /* fppowbf16.vhdl:3971:28  */
  assign n828 = {n826, n827};
  /* fppowbf16.vhdl:3881:10  */
  always @(posedge clk)
    n829 <= sign;
  /* fppowbf16.vhdl:3881:10  */
  always @(posedge clk)
    n830 <= sign_d1;
  /* fppowbf16.vhdl:3881:10  */
  always @(posedge clk)
    n831 <= expx;
  /* fppowbf16.vhdl:3881:10  */
  always @(posedge clk)
    n832 <= expy;
  /* fppowbf16.vhdl:3881:10  */
  always @(posedge clk)
    n833 <= expy_d1;
  /* fppowbf16.vhdl:3881:10  */
  always @(posedge clk)
    n834 <= expy_d2;
  /* fppowbf16.vhdl:3881:10  */
  always @(posedge clk)
    n835 <= expy_d3;
  /* fppowbf16.vhdl:3881:10  */
  always @(posedge clk)
    n836 <= expy_d4;
  /* fppowbf16.vhdl:3881:10  */
  always @(posedge clk)
    n837 <= expy_d5;
  /* fppowbf16.vhdl:3881:10  */
  always @(posedge clk)
    n838 <= expy_d6;
  /* fppowbf16.vhdl:3881:10  */
  always @(posedge clk)
    n839 <= expy_d7;
  /* fppowbf16.vhdl:3881:10  */
  always @(posedge clk)
    n840 <= expy_d8;
  /* fppowbf16.vhdl:3881:10  */
  always @(posedge clk)
    n841 <= expy_d9;
  /* fppowbf16.vhdl:3881:10  */
  always @(posedge clk)
    n842 <= expy_d10;
  /* fppowbf16.vhdl:3881:10  */
  always @(posedge clk)
    n843 <= expy_d11;
  /* fppowbf16.vhdl:3881:10  */
  always @(posedge clk)
    n844 <= expsumpresub;
  /* fppowbf16.vhdl:3881:10  */
  always @(posedge clk)
    n845 <= bias;
  /* fppowbf16.vhdl:3881:10  */
  always @(posedge clk)
    n846 <= bias_d1;
  /* fppowbf16.vhdl:3881:10  */
  always @(posedge clk)
    n847 <= bias_d2;
  /* fppowbf16.vhdl:3881:10  */
  always @(posedge clk)
    n848 <= bias_d3;
  /* fppowbf16.vhdl:3881:10  */
  always @(posedge clk)
    n849 <= bias_d4;
  /* fppowbf16.vhdl:3881:10  */
  always @(posedge clk)
    n850 <= bias_d5;
  /* fppowbf16.vhdl:3881:10  */
  always @(posedge clk)
    n851 <= bias_d6;
  /* fppowbf16.vhdl:3881:10  */
  always @(posedge clk)
    n852 <= bias_d7;
  /* fppowbf16.vhdl:3881:10  */
  always @(posedge clk)
    n853 <= bias_d8;
  /* fppowbf16.vhdl:3881:10  */
  always @(posedge clk)
    n854 <= bias_d9;
  /* fppowbf16.vhdl:3881:10  */
  always @(posedge clk)
    n855 <= bias_d10;
  /* fppowbf16.vhdl:3881:10  */
  always @(posedge clk)
    n856 <= bias_d11;
  /* fppowbf16.vhdl:3881:10  */
  always @(posedge clk)
    n857 <= bias_d12;
  /* fppowbf16.vhdl:3881:10  */
  always @(posedge clk)
    n858 <= sigprod;
  /* fppowbf16.vhdl:3881:10  */
  always @(posedge clk)
    n859 <= exc;
  /* fppowbf16.vhdl:3881:10  */
  always @(posedge clk)
    n860 <= exc_d1;
  /* fppowbf16.vhdl:3881:10  */
  always @(posedge clk)
    n861 <= norm;
  /* fppowbf16.vhdl:3881:10  */
  always @(posedge clk)
    n862 <= norm_d1;
  /* fppowbf16.vhdl:3881:10  */
  always @(posedge clk)
    n863 <= sigprodext;
  /* fppowbf16.vhdl:3881:10  */
  always @(posedge clk)
    n864 <= y;
  /* fppowbf16.vhdl:3881:10  */
  always @(posedge clk)
    n865 <= y_d1;
  /* fppowbf16.vhdl:3881:10  */
  always @(posedge clk)
    n866 <= y_d2;
  /* fppowbf16.vhdl:3881:10  */
  always @(posedge clk)
    n867 <= y_d3;
  /* fppowbf16.vhdl:3881:10  */
  always @(posedge clk)
    n868 <= y_d4;
  /* fppowbf16.vhdl:3881:10  */
  always @(posedge clk)
    n869 <= y_d5;
  /* fppowbf16.vhdl:3881:10  */
  always @(posedge clk)
    n870 <= y_d6;
  /* fppowbf16.vhdl:3881:10  */
  always @(posedge clk)
    n871 <= y_d7;
  /* fppowbf16.vhdl:3881:10  */
  always @(posedge clk)
    n872 <= y_d8;
  /* fppowbf16.vhdl:3881:10  */
  always @(posedge clk)
    n873 <= y_d9;
  /* fppowbf16.vhdl:3881:10  */
  always @(posedge clk)
    n874 <= y_d10;
endmodule

module fplogiterative_8_17_0_500_freq500_uid9
  (input  clk,
   input  [27:0] x,
   output [27:0] r);
  wire [2:0] xexnsgn;
  wire [2:0] xexnsgn_d1;
  wire [2:0] xexnsgn_d2;
  wire [2:0] xexnsgn_d3;
  wire [2:0] xexnsgn_d4;
  wire [2:0] xexnsgn_d5;
  wire [2:0] xexnsgn_d6;
  wire [2:0] xexnsgn_d7;
  wire [2:0] xexnsgn_d8;
  wire [2:0] xexnsgn_d9;
  wire [2:0] xexnsgn_d10;
  wire [2:0] xexnsgn_d11;
  wire firstbit;
  wire [18:0] y0;
  wire [18:0] y0_d1;
  wire [16:0] y0h;
  wire sr;
  wire sr_d1;
  wire sr_d2;
  wire sr_d3;
  wire sr_d4;
  wire sr_d5;
  wire sr_d6;
  wire sr_d7;
  wire sr_d8;
  wire sr_d9;
  wire sr_d10;
  wire sr_d11;
  wire [9:0] absz0;
  wire [7:0] e;
  wire [7:0] abse;
  wire eeqzero;
  wire eeqzero_d1;
  wire eeqzero_d2;
  wire eeqzero_d3;
  wire eeqzero_d4;
  wire [4:0] lzo;
  wire [4:0] lzo_d1;
  wire [4:0] lzo_d2;
  wire [4:0] lzo_d3;
  wire [4:0] pfinal_s;
  wire [4:0] pfinal_s_d1;
  wire [4:0] pfinal_s_d2;
  wire [4:0] pfinal_s_d3;
  wire [5:0] shiftval;
  wire [3:0] shiftvalinl;
  wire [3:0] shiftvalinr;
  wire dorr;
  wire dorr_d1;
  wire dorr_d2;
  wire \small ;
  wire small_d1;
  wire small_d2;
  wire small_d3;
  wire small_d4;
  wire small_d5;
  wire small_d6;
  wire small_d7;
  wire [19:0] small_absz0_normd_full;
  wire [9:0] small_absz0_normd;
  wire [9:0] small_absz0_normd_d1;
  wire [6:0] a0;
  wire [7:0] inva0;
  wire [7:0] inva0_d1;
  wire [7:0] inva0_copy16;
  wire [26:0] p0;
  wire [19:0] z1;
  wire [4:0] a1;
  wire [4:0] a1_d1;
  wire [14:0] b1;
  wire [19:0] zm1;
  wire [19:0] zm1_d1;
  wire [24:0] p1;
  wire [25:0] y1;
  wire [20:0] eiy1;
  wire [20:0] addxiter1;
  wire [20:0] eiypb1;
  wire [20:0] pp1;
  wire [20:0] z2;
  wire [20:0] zfinal;
  wire [20:0] zfinal_d1;
  wire [20:0] zfinal_d2;
  wire [13:0] squarerin;
  wire [27:0] z2o2_full;
  wire [27:0] z2o2_full_dummy;
  wire [10:0] z2o2_normal;
  wire [20:0] addfinallog1py;
  wire [20:0] log1p_normal;
  wire [29:0] l0;
  wire [29:0] l0_copy28;
  wire [29:0] s1;
  wire [24:0] l1;
  wire [24:0] l1_copy31;
  wire [29:0] sopx1;
  wire [29:0] s2;
  wire [29:0] almostlog;
  wire [29:0] adderlogf_normaly;
  wire [29:0] logf_normal;
  wire [28:0] abselog2;
  wire [37:0] abselog2_pad;
  wire [37:0] logf_normal_pad;
  wire [37:0] lnaddx;
  wire [37:0] lnaddy;
  wire [37:0] log_normal;
  wire [29:0] log_normal_normd;
  wire [4:0] e_normal;
  wire [13:0] z2o2_small_bs;
  wire [26:0] z2o2_small_s;
  wire [22:0] z2o2_small;
  wire [22:0] z_small;
  wire [22:0] log_smally;
  wire nsrcin;
  wire [22:0] log_small;
  wire [1:0] e0_sub;
  wire ufl;
  wire ufl_d1;
  wire ufl_d2;
  wire ufl_d3;
  wire ufl_d4;
  wire ufl_d5;
  wire ufl_d6;
  wire ufl_d7;
  wire ufl_d8;
  wire ufl_d9;
  wire ufl_d10;
  wire ufl_d11;
  wire [7:0] e_small;
  wire [7:0] e_small_d1;
  wire [7:0] e_small_d2;
  wire [7:0] e_small_d3;
  wire [7:0] e_small_d4;
  wire [20:0] log_small_normd;
  wire [20:0] log_small_normd_d1;
  wire [20:0] log_small_normd_d2;
  wire [20:0] log_small_normd_d3;
  wire [20:0] log_small_normd_d4;
  wire [20:0] log_small_normd_d5;
  wire [7:0] e0offset;
  wire [7:0] e0offset_d1;
  wire [7:0] e0offset_d2;
  wire [7:0] e0offset_d3;
  wire [7:0] e0offset_d4;
  wire [7:0] e0offset_d5;
  wire [7:0] e0offset_d6;
  wire [7:0] e0offset_d7;
  wire [7:0] e0offset_d8;
  wire [7:0] e0offset_d9;
  wire [7:0] e0offset_d10;
  wire [7:0] er;
  wire [7:0] er_d1;
  wire [20:0] log_g;
  wire round;
  wire [24:0] frax;
  wire [24:0] fray;
  wire [24:0] efr;
  wire [2:0] rexn;
  wire [2:0] n356;
  wire n357;
  wire [16:0] n358;
  wire [17:0] n360;
  wire [18:0] n362;
  wire n363;
  wire [18:0] n364;
  wire [16:0] n365;
  wire [18:0] n367;
  wire [16:0] n368;
  wire [7:0] n370;
  wire n372;
  wire n373;
  wire n374;
  wire n375;
  wire [9:0] n376;
  wire n377;
  wire [9:0] n378;
  wire [9:0] n379;
  wire [9:0] n381;
  wire [7:0] n382;
  wire n383;
  wire [7:0] n385;
  wire [7:0] n386;
  wire [7:0] n388;
  wire [7:0] n389;
  wire n392;
  wire n393;
  wire [4:0] lzoc1_n395;
  wire [5:0] n400;
  wire [5:0] n402;
  wire [5:0] n403;
  wire [3:0] n404;
  wire [3:0] n405;
  wire n406;
  wire n407;
  wire n408;
  wire [19:0] small_lshift_n409;
  wire [9:0] n412;
  wire [6:0] n413;
  wire [7:0] inva0table_n414;
  wire [26:0] n417;
  wire [26:0] n418;
  wire [26:0] n419;
  wire [19:0] n420;
  wire [4:0] n421;
  wire [14:0] n422;
  wire [24:0] n423;
  wire [24:0] n424;
  wire [24:0] n425;
  wire [25:0] n427;
  wire [20:0] n428;
  wire n429;
  wire [20:0] n430;
  wire [19:0] n431;
  wire [20:0] n433;
  wire [15:0] n435;
  wire [20:0] n437;
  localparam n438 = 1'b0;
  wire [20:0] additer1_1_n439;
  wire [19:0] n442;
  wire [19:0] n443;
  wire [20:0] n445;
  localparam n446 = 1'b1;
  wire [20:0] additer2_1_n447;
  wire [13:0] n450;
  wire [13:0] n451;
  wire [13:0] n453;
  wire [27:0] n454;
  wire [27:0] n455;
  wire [27:0] n456;
  wire [10:0] n457;
  wire [10:0] n458;
  wire [20:0] n460;
  localparam n461 = 1'b1;
  wire [20:0] addfinallog1p_normaladder_n462;
  wire [29:0] logtable0_n465;
  wire [24:0] logtable1_n468;
  wire [29:0] n472;
  localparam n473 = 1'b0;
  wire [29:0] adders1_n474;
  wire [29:0] n478;
  localparam n479 = 1'b0;
  wire [29:0] adderlogf_normal_n480;
  wire [28:0] mullog2_n483;
  wire [37:0] n487;
  wire n488;
  wire n489;
  wire n490;
  wire n491;
  wire n492;
  wire n493;
  wire n494;
  wire n495;
  wire [3:0] n496;
  wire [3:0] n497;
  wire [7:0] n498;
  wire [37:0] n499;
  wire n500;
  wire [37:0] n501;
  wire [37:0] n502;
  wire [37:0] lnadder_n503;
  wire [4:0] final_norm_n506;
  wire [29:0] final_norm_n507;
  wire [13:0] n512;
  wire [26:0] ao_rshift_n513;
  wire [13:0] n516;
  wire [22:0] n518;
  wire [22:0] n520;
  wire [22:0] n521;
  wire [22:0] n522;
  wire n523;
  wire [22:0] log_small_adder_n524;
  wire n528;
  wire [1:0] n529;
  wire [1:0] n531;
  wire n533;
  wire [1:0] n534;
  wire [7:0] n538;
  wire [7:0] n540;
  wire [7:0] n541;
  wire [20:0] n542;
  wire n543;
  wire [20:0] n544;
  wire [20:0] n545;
  wire n546;
  wire [20:0] n547;
  wire [20:0] n548;
  wire [7:0] n550;
  wire [7:0] n552;
  wire [7:0] n553;
  wire [19:0] n554;
  wire [20:0] n556;
  wire [20:0] n557;
  wire [20:0] n558;
  wire n559;
  wire [16:0] n560;
  wire [24:0] n561;
  wire [24:0] n563;
  localparam n564 = 1'b0;
  wire [24:0] finalroundadder_n565;
  wire n569;
  wire n570;
  wire n571;
  wire n572;
  wire n573;
  wire n574;
  wire n575;
  wire n576;
  wire n577;
  wire [2:0] n578;
  wire [1:0] n580;
  wire n582;
  wire [2:0] n583;
  wire [1:0] n585;
  wire n587;
  wire [2:0] n588;
  wire [2:0] n590;
  wire n591;
  wire n592;
  wire n593;
  wire n594;
  wire n595;
  wire n596;
  wire n597;
  wire n598;
  wire n599;
  wire n600;
  wire [2:0] n601;
  wire [2:0] n603;
  wire [27:0] n604;
  reg [2:0] n605;
  reg [2:0] n606;
  reg [2:0] n607;
  reg [2:0] n608;
  reg [2:0] n609;
  reg [2:0] n610;
  reg [2:0] n611;
  reg [2:0] n612;
  reg [2:0] n613;
  reg [2:0] n614;
  reg [2:0] n615;
  reg [18:0] n616;
  reg n617;
  reg n618;
  reg n619;
  reg n620;
  reg n621;
  reg n622;
  reg n623;
  reg n624;
  reg n625;
  reg n626;
  reg n627;
  reg n628;
  reg n629;
  reg n630;
  reg n631;
  reg [4:0] n632;
  reg [4:0] n633;
  reg [4:0] n634;
  reg [4:0] n635;
  reg [4:0] n636;
  reg [4:0] n637;
  reg n638;
  reg n639;
  reg n640;
  reg n641;
  reg n642;
  reg n643;
  reg n644;
  reg n645;
  reg n646;
  reg [9:0] n647;
  reg [7:0] n648;
  reg [4:0] n649;
  reg [19:0] n650;
  reg [20:0] n651;
  reg [20:0] n652;
  reg n653;
  reg n654;
  reg n655;
  reg n656;
  reg n657;
  reg n658;
  reg n659;
  reg n660;
  reg n661;
  reg n662;
  reg n663;
  reg [7:0] n664;
  reg [7:0] n665;
  reg [7:0] n666;
  reg [7:0] n667;
  reg [20:0] n668;
  reg [20:0] n669;
  reg [20:0] n670;
  reg [20:0] n671;
  reg [20:0] n672;
  reg [7:0] n673;
  reg [7:0] n674;
  reg [7:0] n675;
  reg [7:0] n676;
  reg [7:0] n677;
  reg [7:0] n678;
  reg [7:0] n679;
  reg [7:0] n680;
  reg [7:0] n681;
  reg [7:0] n682;
  reg [7:0] n683;
  assign r = n604; //(module output)
  /* fppowbf16.vhdl:3234:8  */
  assign xexnsgn = n356; // (signal)
  /* fppowbf16.vhdl:3234:17  */
  assign xexnsgn_d1 = n605; // (signal)
  /* fppowbf16.vhdl:3234:29  */
  assign xexnsgn_d2 = n606; // (signal)
  /* fppowbf16.vhdl:3234:41  */
  assign xexnsgn_d3 = n607; // (signal)
  /* fppowbf16.vhdl:3234:53  */
  assign xexnsgn_d4 = n608; // (signal)
  /* fppowbf16.vhdl:3234:65  */
  assign xexnsgn_d5 = n609; // (signal)
  /* fppowbf16.vhdl:3234:77  */
  assign xexnsgn_d6 = n610; // (signal)
  /* fppowbf16.vhdl:3234:89  */
  assign xexnsgn_d7 = n611; // (signal)
  /* fppowbf16.vhdl:3234:101  */
  assign xexnsgn_d8 = n612; // (signal)
  /* fppowbf16.vhdl:3234:113  */
  assign xexnsgn_d9 = n613; // (signal)
  /* fppowbf16.vhdl:3234:125  */
  assign xexnsgn_d10 = n614; // (signal)
  /* fppowbf16.vhdl:3234:138  */
  assign xexnsgn_d11 = n615; // (signal)
  /* fppowbf16.vhdl:3236:8  */
  assign firstbit = n357; // (signal)
  /* fppowbf16.vhdl:3238:8  */
  assign y0 = n364; // (signal)
  /* fppowbf16.vhdl:3238:12  */
  assign y0_d1 = n616; // (signal)
  /* fppowbf16.vhdl:3240:8  */
  assign y0h = n368; // (signal)
  /* fppowbf16.vhdl:3242:8  */
  assign sr = n373; // (signal)
  /* fppowbf16.vhdl:3242:12  */
  assign sr_d1 = n617; // (signal)
  /* fppowbf16.vhdl:3242:19  */
  assign sr_d2 = n618; // (signal)
  /* fppowbf16.vhdl:3242:26  */
  assign sr_d3 = n619; // (signal)
  /* fppowbf16.vhdl:3242:33  */
  assign sr_d4 = n620; // (signal)
  /* fppowbf16.vhdl:3242:40  */
  assign sr_d5 = n621; // (signal)
  /* fppowbf16.vhdl:3242:47  */
  assign sr_d6 = n622; // (signal)
  /* fppowbf16.vhdl:3242:54  */
  assign sr_d7 = n623; // (signal)
  /* fppowbf16.vhdl:3242:61  */
  assign sr_d8 = n624; // (signal)
  /* fppowbf16.vhdl:3242:68  */
  assign sr_d9 = n625; // (signal)
  /* fppowbf16.vhdl:3242:75  */
  assign sr_d10 = n626; // (signal)
  /* fppowbf16.vhdl:3242:83  */
  assign sr_d11 = n627; // (signal)
  /* fppowbf16.vhdl:3244:8  */
  assign absz0 = n378; // (signal)
  /* fppowbf16.vhdl:3246:8  */
  assign e = n386; // (signal)
  /* fppowbf16.vhdl:3248:8  */
  assign abse = n389; // (signal)
  /* fppowbf16.vhdl:3250:8  */
  assign eeqzero = n393; // (signal)
  /* fppowbf16.vhdl:3250:17  */
  assign eeqzero_d1 = n628; // (signal)
  /* fppowbf16.vhdl:3250:29  */
  assign eeqzero_d2 = n629; // (signal)
  /* fppowbf16.vhdl:3250:41  */
  assign eeqzero_d3 = n630; // (signal)
  /* fppowbf16.vhdl:3250:53  */
  assign eeqzero_d4 = n631; // (signal)
  /* fppowbf16.vhdl:3252:8  */
  assign lzo = lzoc1_n395; // (signal)
  /* fppowbf16.vhdl:3252:13  */
  assign lzo_d1 = n632; // (signal)
  /* fppowbf16.vhdl:3252:21  */
  assign lzo_d2 = n633; // (signal)
  /* fppowbf16.vhdl:3252:29  */
  assign lzo_d3 = n634; // (signal)
  /* fppowbf16.vhdl:3254:8  */
  assign pfinal_s = 5'b01001; // (signal)
  /* fppowbf16.vhdl:3254:18  */
  assign pfinal_s_d1 = n635; // (signal)
  /* fppowbf16.vhdl:3254:31  */
  assign pfinal_s_d2 = n636; // (signal)
  /* fppowbf16.vhdl:3254:44  */
  assign pfinal_s_d3 = n637; // (signal)
  /* fppowbf16.vhdl:3256:8  */
  assign shiftval = n403; // (signal)
  /* fppowbf16.vhdl:3258:8  */
  assign shiftvalinl = n404; // (signal)
  /* fppowbf16.vhdl:3260:8  */
  assign shiftvalinr = n405; // (signal)
  /* fppowbf16.vhdl:3262:8  */
  assign dorr = n406; // (signal)
  /* fppowbf16.vhdl:3262:14  */
  assign dorr_d1 = n638; // (signal)
  /* fppowbf16.vhdl:3262:23  */
  assign dorr_d2 = n639; // (signal)
  /* fppowbf16.vhdl:3264:8  */
  assign \small  = n408; // (signal)
  /* fppowbf16.vhdl:3264:15  */
  assign small_d1 = n640; // (signal)
  /* fppowbf16.vhdl:3264:25  */
  assign small_d2 = n641; // (signal)
  /* fppowbf16.vhdl:3264:35  */
  assign small_d3 = n642; // (signal)
  /* fppowbf16.vhdl:3264:45  */
  assign small_d4 = n643; // (signal)
  /* fppowbf16.vhdl:3264:55  */
  assign small_d5 = n644; // (signal)
  /* fppowbf16.vhdl:3264:65  */
  assign small_d6 = n645; // (signal)
  /* fppowbf16.vhdl:3264:75  */
  assign small_d7 = n646; // (signal)
  /* fppowbf16.vhdl:3266:8  */
  assign small_absz0_normd_full = small_lshift_n409; // (signal)
  /* fppowbf16.vhdl:3268:8  */
  assign small_absz0_normd = n412; // (signal)
  /* fppowbf16.vhdl:3268:27  */
  assign small_absz0_normd_d1 = n647; // (signal)
  /* fppowbf16.vhdl:3270:8  */
  assign a0 = n413; // (signal)
  /* fppowbf16.vhdl:3272:8  */
  assign inva0 = inva0_copy16; // (signal)
  /* fppowbf16.vhdl:3272:15  */
  assign inva0_d1 = n648; // (signal)
  /* fppowbf16.vhdl:3274:8  */
  assign inva0_copy16 = inva0table_n414; // (signal)
  /* fppowbf16.vhdl:3276:8  */
  assign p0 = n419; // (signal)
  /* fppowbf16.vhdl:3278:8  */
  assign z1 = n420; // (signal)
  /* fppowbf16.vhdl:3280:8  */
  assign a1 = n421; // (signal)
  /* fppowbf16.vhdl:3280:12  */
  assign a1_d1 = n649; // (signal)
  /* fppowbf16.vhdl:3282:8  */
  assign b1 = n422; // (signal)
  /* fppowbf16.vhdl:3284:8  */
  assign zm1 = z1; // (signal)
  /* fppowbf16.vhdl:3284:13  */
  assign zm1_d1 = n650; // (signal)
  /* fppowbf16.vhdl:3286:8  */
  assign p1 = n425; // (signal)
  /* fppowbf16.vhdl:3288:8  */
  assign y1 = n427; // (signal)
  /* fppowbf16.vhdl:3290:8  */
  assign eiy1 = n430; // (signal)
  /* fppowbf16.vhdl:3292:8  */
  assign addxiter1 = n437; // (signal)
  /* fppowbf16.vhdl:3294:8  */
  assign eiypb1 = additer1_1_n439; // (signal)
  /* fppowbf16.vhdl:3296:8  */
  assign pp1 = n445; // (signal)
  /* fppowbf16.vhdl:3298:8  */
  assign z2 = additer2_1_n447; // (signal)
  /* fppowbf16.vhdl:3300:8  */
  assign zfinal = z2; // (signal)
  /* fppowbf16.vhdl:3300:16  */
  assign zfinal_d1 = n651; // (signal)
  /* fppowbf16.vhdl:3300:27  */
  assign zfinal_d2 = n652; // (signal)
  /* fppowbf16.vhdl:3302:8  */
  assign squarerin = n451; // (signal)
  /* fppowbf16.vhdl:3304:8  */
  assign z2o2_full = n456; // (signal)
  /* fppowbf16.vhdl:3306:8  */
  assign z2o2_full_dummy = z2o2_full; // (signal)
  /* fppowbf16.vhdl:3308:8  */
  assign z2o2_normal = n457; // (signal)
  /* fppowbf16.vhdl:3310:8  */
  assign addfinallog1py = n460; // (signal)
  /* fppowbf16.vhdl:3312:8  */
  assign log1p_normal = addfinallog1p_normaladder_n462; // (signal)
  /* fppowbf16.vhdl:3314:8  */
  assign l0 = l0_copy28; // (signal)
  /* fppowbf16.vhdl:3316:8  */
  assign l0_copy28 = logtable0_n465; // (signal)
  /* fppowbf16.vhdl:3318:8  */
  assign s1 = l0; // (signal)
  /* fppowbf16.vhdl:3320:8  */
  assign l1 = l1_copy31; // (signal)
  /* fppowbf16.vhdl:3322:8  */
  assign l1_copy31 = logtable1_n468; // (signal)
  /* fppowbf16.vhdl:3324:8  */
  assign sopx1 = n472; // (signal)
  /* fppowbf16.vhdl:3326:8  */
  assign s2 = adders1_n474; // (signal)
  /* fppowbf16.vhdl:3328:8  */
  assign almostlog = s2; // (signal)
  /* fppowbf16.vhdl:3330:8  */
  assign adderlogf_normaly = n478; // (signal)
  /* fppowbf16.vhdl:3332:8  */
  assign logf_normal = adderlogf_normal_n480; // (signal)
  /* fppowbf16.vhdl:3334:8  */
  assign abselog2 = mullog2_n483; // (signal)
  /* fppowbf16.vhdl:3336:8  */
  assign abselog2_pad = n487; // (signal)
  /* fppowbf16.vhdl:3338:8  */
  assign logf_normal_pad = n499; // (signal)
  /* fppowbf16.vhdl:3340:8  */
  assign lnaddx = abselog2_pad; // (signal)
  /* fppowbf16.vhdl:3342:8  */
  assign lnaddy = n501; // (signal)
  /* fppowbf16.vhdl:3344:8  */
  assign log_normal = lnadder_n503; // (signal)
  /* fppowbf16.vhdl:3346:8  */
  assign log_normal_normd = final_norm_n507; // (signal)
  /* fppowbf16.vhdl:3348:8  */
  assign e_normal = final_norm_n506; // (signal)
  /* fppowbf16.vhdl:3350:8  */
  assign z2o2_small_bs = n512; // (signal)
  /* fppowbf16.vhdl:3352:8  */
  assign z2o2_small_s = ao_rshift_n513; // (signal)
  /* fppowbf16.vhdl:3354:8  */
  assign z2o2_small = n518; // (signal)
  /* fppowbf16.vhdl:3356:8  */
  assign z_small = n520; // (signal)
  /* fppowbf16.vhdl:3358:8  */
  assign log_smally = n521; // (signal)
  /* fppowbf16.vhdl:3360:8  */
  assign nsrcin = n523; // (signal)
  /* fppowbf16.vhdl:3362:8  */
  assign log_small = log_small_adder_n524; // (signal)
  /* fppowbf16.vhdl:3364:8  */
  assign e0_sub = n529; // (signal)
  /* fppowbf16.vhdl:3366:8  */
  assign ufl = 1'b0; // (signal)
  /* fppowbf16.vhdl:3366:13  */
  assign ufl_d1 = n653; // (signal)
  /* fppowbf16.vhdl:3366:21  */
  assign ufl_d2 = n654; // (signal)
  /* fppowbf16.vhdl:3366:29  */
  assign ufl_d3 = n655; // (signal)
  /* fppowbf16.vhdl:3366:37  */
  assign ufl_d4 = n656; // (signal)
  /* fppowbf16.vhdl:3366:45  */
  assign ufl_d5 = n657; // (signal)
  /* fppowbf16.vhdl:3366:53  */
  assign ufl_d6 = n658; // (signal)
  /* fppowbf16.vhdl:3366:61  */
  assign ufl_d7 = n659; // (signal)
  /* fppowbf16.vhdl:3366:69  */
  assign ufl_d8 = n660; // (signal)
  /* fppowbf16.vhdl:3366:77  */
  assign ufl_d9 = n661; // (signal)
  /* fppowbf16.vhdl:3366:85  */
  assign ufl_d10 = n662; // (signal)
  /* fppowbf16.vhdl:3366:94  */
  assign ufl_d11 = n663; // (signal)
  /* fppowbf16.vhdl:3368:8  */
  assign e_small = n541; // (signal)
  /* fppowbf16.vhdl:3368:17  */
  assign e_small_d1 = n664; // (signal)
  /* fppowbf16.vhdl:3368:29  */
  assign e_small_d2 = n665; // (signal)
  /* fppowbf16.vhdl:3368:41  */
  assign e_small_d3 = n666; // (signal)
  /* fppowbf16.vhdl:3368:53  */
  assign e_small_d4 = n667; // (signal)
  /* fppowbf16.vhdl:3370:8  */
  assign log_small_normd = n544; // (signal)
  /* fppowbf16.vhdl:3370:25  */
  assign log_small_normd_d1 = n668; // (signal)
  /* fppowbf16.vhdl:3370:45  */
  assign log_small_normd_d2 = n669; // (signal)
  /* fppowbf16.vhdl:3370:65  */
  assign log_small_normd_d3 = n670; // (signal)
  /* fppowbf16.vhdl:3370:85  */
  assign log_small_normd_d4 = n671; // (signal)
  /* fppowbf16.vhdl:3370:105  */
  assign log_small_normd_d5 = n672; // (signal)
  /* fppowbf16.vhdl:3372:8  */
  assign e0offset = 8'b10000110; // (signal)
  /* fppowbf16.vhdl:3372:18  */
  assign e0offset_d1 = n673; // (signal)
  /* fppowbf16.vhdl:3372:31  */
  assign e0offset_d2 = n674; // (signal)
  /* fppowbf16.vhdl:3372:44  */
  assign e0offset_d3 = n675; // (signal)
  /* fppowbf16.vhdl:3372:57  */
  assign e0offset_d4 = n676; // (signal)
  /* fppowbf16.vhdl:3372:70  */
  assign e0offset_d5 = n677; // (signal)
  /* fppowbf16.vhdl:3372:83  */
  assign e0offset_d6 = n678; // (signal)
  /* fppowbf16.vhdl:3372:96  */
  assign e0offset_d7 = n679; // (signal)
  /* fppowbf16.vhdl:3372:109  */
  assign e0offset_d8 = n680; // (signal)
  /* fppowbf16.vhdl:3372:122  */
  assign e0offset_d9 = n681; // (signal)
  /* fppowbf16.vhdl:3372:135  */
  assign e0offset_d10 = n682; // (signal)
  /* fppowbf16.vhdl:3374:8  */
  assign er = n550; // (signal)
  /* fppowbf16.vhdl:3374:12  */
  assign er_d1 = n683; // (signal)
  /* fppowbf16.vhdl:3376:8  */
  assign log_g = n557; // (signal)
  /* fppowbf16.vhdl:3378:8  */
  assign round = n559; // (signal)
  /* fppowbf16.vhdl:3380:8  */
  assign frax = n561; // (signal)
  /* fppowbf16.vhdl:3382:8  */
  assign fray = n563; // (signal)
  /* fppowbf16.vhdl:3384:8  */
  assign efr = finalroundadder_n565; // (signal)
  /* fppowbf16.vhdl:3386:8  */
  assign rexn = n578; // (signal)
  /* fppowbf16.vhdl:3480:17  */
  assign n356 = x[27:25]; // extract
  /* fppowbf16.vhdl:3481:18  */
  assign n357 = x[16]; // extract
  /* fppowbf16.vhdl:3482:17  */
  assign n358 = x[16:0]; // extract
  /* fppowbf16.vhdl:3482:14  */
  assign n360 = {1'b1, n358};
  /* fppowbf16.vhdl:3482:33  */
  assign n362 = {n360, 1'b0};
  /* fppowbf16.vhdl:3482:53  */
  assign n363 = ~firstbit;
  /* fppowbf16.vhdl:3482:39  */
  assign n364 = n363 ? n362 : n367;
  /* fppowbf16.vhdl:3482:72  */
  assign n365 = x[16:0]; // extract
  /* fppowbf16.vhdl:3482:69  */
  assign n367 = {2'b01, n365};
  /* fppowbf16.vhdl:3483:13  */
  assign n368 = y0[17:1]; // extract
  /* fppowbf16.vhdl:3485:24  */
  assign n370 = x[24:17]; // extract
  /* fppowbf16.vhdl:3485:44  */
  assign n372 = n370 == 8'b01111111;
  /* fppowbf16.vhdl:3485:16  */
  assign n373 = n372 ? 1'b0 : n375;
  /* fppowbf16.vhdl:3486:16  */
  assign n374 = x[24]; // extract
  /* fppowbf16.vhdl:3486:11  */
  assign n375 = ~n374;
  /* fppowbf16.vhdl:3487:17  */
  assign n376 = y0[9:0]; // extract
  /* fppowbf16.vhdl:3487:57  */
  assign n377 = ~sr;
  /* fppowbf16.vhdl:3487:49  */
  assign n378 = n377 ? n376 : n381;
  /* fppowbf16.vhdl:3488:49  */
  assign n379 = y0[9:0]; // extract
  /* fppowbf16.vhdl:3488:45  */
  assign n381 = 10'b0000000000 - n379;
  /* fppowbf16.vhdl:3489:11  */
  assign n382 = x[24:17]; // extract
  /* fppowbf16.vhdl:3489:67  */
  assign n383 = ~firstbit;
  /* fppowbf16.vhdl:3489:64  */
  assign n385 = {7'b0111111, n383};
  /* fppowbf16.vhdl:3489:32  */
  assign n386 = n382 - n385;
  /* fppowbf16.vhdl:3490:36  */
  assign n388 = 8'b00000000 - e;
  /* fppowbf16.vhdl:3490:43  */
  assign n389 = sr ? n388 : e;
  /* fppowbf16.vhdl:3491:25  */
  assign n392 = e == 8'b00000000;
  /* fppowbf16.vhdl:3491:19  */
  assign n393 = n392 ? 1'b1 : 1'b0;
  /* fppowbf16.vhdl:3492:4  */
  lzoc_17_freq500_uid11 lzoc1 (
    .clk(clk),
    .i(y0h),
    .ozb(firstbit),
    .o(lzoc1_n395));
  /* fppowbf16.vhdl:3498:21  */
  assign n400 = {1'b0, lzo};
  /* fppowbf16.vhdl:3498:35  */
  assign n402 = {1'b0, pfinal_s_d3};
  /* fppowbf16.vhdl:3498:28  */
  assign n403 = n400 - n402;
  /* fppowbf16.vhdl:3499:27  */
  assign n404 = shiftval[3:0]; // extract
  /* fppowbf16.vhdl:3500:27  */
  assign n405 = shiftval[3:0]; // extract
  /* fppowbf16.vhdl:3501:20  */
  assign n406 = shiftval[5]; // extract
  /* fppowbf16.vhdl:3502:28  */
  assign n407 = ~dorr_d1;
  /* fppowbf16.vhdl:3502:24  */
  assign n408 = eeqzero_d4 & n407;
  /* fppowbf16.vhdl:3504:4  */
  leftshifter10_by_max_10_freq500_uid13 small_lshift (
    .clk(clk),
    .x(absz0),
    .s(shiftvalinl),
    .r(small_lshift_n409));
  /* fppowbf16.vhdl:3509:47  */
  assign n412 = small_absz0_normd_full[9:0]; // extract
  /* fppowbf16.vhdl:3511:11  */
  assign n413 = x[16:10]; // extract
  /* fppowbf16.vhdl:3513:4  */
  inva0table_freq500_uid15 inva0table (
    .x(a0),
    .y(inva0table_n414));
  /* fppowbf16.vhdl:3517:19  */
  assign n417 = {19'b0, inva0_d1};  //  uext
  /* fppowbf16.vhdl:3517:19  */
  assign n418 = {8'b0, y0_d1};  //  uext
  /* fppowbf16.vhdl:3517:19  */
  assign n419 = n417 * n418; // umul
  /* fppowbf16.vhdl:3519:12  */
  assign n420 = p0[19:0]; // extract
  /* fppowbf16.vhdl:3521:12  */
  assign n421 = z1[19:15]; // extract
  /* fppowbf16.vhdl:3522:12  */
  assign n422 = z1[14:0]; // extract
  /* fppowbf16.vhdl:3524:15  */
  assign n423 = {20'b0, a1_d1};  //  uext
  /* fppowbf16.vhdl:3524:15  */
  assign n424 = {5'b0, zm1_d1};  //  uext
  /* fppowbf16.vhdl:3524:15  */
  assign n425 = n423 * n424; // umul
  /* fppowbf16.vhdl:3525:36  */
  assign n427 = {6'b100000, z1};
  /* fppowbf16.vhdl:3526:14  */
  assign n428 = y1[25:5]; // extract
  /* fppowbf16.vhdl:3526:36  */
  assign n429 = a1[4]; // extract
  /* fppowbf16.vhdl:3526:29  */
  assign n430 = n429 ? n428 : n433;
  /* fppowbf16.vhdl:3527:20  */
  assign n431 = y1[25:6]; // extract
  /* fppowbf16.vhdl:3527:16  */
  assign n433 = {1'b0, n431};
  /* fppowbf16.vhdl:3528:21  */
  assign n435 = {1'b0, b1};
  /* fppowbf16.vhdl:3528:26  */
  assign n437 = {n435, 5'b00000};
  /* fppowbf16.vhdl:3529:4  */
  intadder_21_freq500_uid19 additer1_1 (
    .clk(clk),
    .x(addxiter1),
    .y(eiy1),
    .cin(n438),
    .r(additer1_1_n439));
  /* fppowbf16.vhdl:3535:39  */
  assign n442 = p1[24:5]; // extract
  /* fppowbf16.vhdl:3535:33  */
  assign n443 = ~n442;
  /* fppowbf16.vhdl:3535:31  */
  assign n445 = {1'b1, n443};
  /* fppowbf16.vhdl:3536:4  */
  intadder_21_freq500_uid22 additer2_1 (
    .clk(clk),
    .x(eiypb1),
    .y(pp1),
    .cin(n446),
    .r(additer2_1_n447));
  /* fppowbf16.vhdl:3543:26  */
  assign n450 = zfinal_d2[20:7]; // extract
  /* fppowbf16.vhdl:3543:54  */
  assign n451 = dorr_d2 ? n450 : n453;
  /* fppowbf16.vhdl:3544:48  */
  assign n453 = {small_absz0_normd_d1, 4'b0000};
  /* fppowbf16.vhdl:3545:26  */
  assign n454 = {14'b0, squarerin};  //  uext
  /* fppowbf16.vhdl:3545:26  */
  assign n455 = {14'b0, squarerin};  //  uext
  /* fppowbf16.vhdl:3545:26  */
  assign n456 = n454 * n455; // umul
  /* fppowbf16.vhdl:3547:35  */
  assign n457 = z2o2_full_dummy[27:17]; // extract
  /* fppowbf16.vhdl:3548:50  */
  assign n458 = ~z2o2_normal;
  /* fppowbf16.vhdl:3548:48  */
  assign n460 = {10'b1111111111, n458};
  /* fppowbf16.vhdl:3549:4  */
  intadder_21_freq500_uid25 addfinallog1p_normaladder (
    .clk(clk),
    .x(zfinal),
    .y(addfinallog1py),
    .cin(n461),
    .r(addfinallog1p_normaladder_n462));
  /* fppowbf16.vhdl:3557:4  */
  logtable0_freq500_uid27 logtable0 (
    .x(a0),
    .y(logtable0_n465));
  /* fppowbf16.vhdl:3562:4  */
  logtable1_freq500_uid30 logtable1 (
    .x(a1),
    .y(logtable1_n468));
  /* fppowbf16.vhdl:3566:36  */
  assign n472 = {5'b00000, l1};
  /* fppowbf16.vhdl:3567:4  */
  intadder_30_freq500_uid34 adders1 (
    .clk(clk),
    .x(s1),
    .y(sopx1),
    .cin(n473),
    .r(adders1_n474));
  /* fppowbf16.vhdl:3574:62  */
  assign n478 = {9'b000000000, log1p_normal};
  /* fppowbf16.vhdl:3575:4  */
  intadder_30_freq500_uid37 adderlogf_normal (
    .clk(clk),
    .x(almostlog),
    .y(adderlogf_normaly),
    .cin(n479),
    .r(adderlogf_normal_n480));
  /* fppowbf16.vhdl:3581:4  */
  fixrealkcm_freq500_uid39 mullog2 (
    .clk(clk),
    .x(abse),
    .r(mullog2_n483));
  /* fppowbf16.vhdl:3585:31  */
  assign n487 = {abselog2, 9'b000000000};
  /* fppowbf16.vhdl:3586:53  */
  assign n488 = logf_normal[29]; // extract
  /* fppowbf16.vhdl:3586:53  */
  assign n489 = logf_normal[29]; // extract
  /* fppowbf16.vhdl:3586:53  */
  assign n490 = logf_normal[29]; // extract
  /* fppowbf16.vhdl:3586:53  */
  assign n491 = logf_normal[29]; // extract
  /* fppowbf16.vhdl:3586:53  */
  assign n492 = logf_normal[29]; // extract
  /* fppowbf16.vhdl:3586:53  */
  assign n493 = logf_normal[29]; // extract
  /* fppowbf16.vhdl:3586:53  */
  assign n494 = logf_normal[29]; // extract
  /* fppowbf16.vhdl:3586:53  */
  assign n495 = logf_normal[29]; // extract
  assign n496 = {n495, n494, n493, n492};
  assign n497 = {n491, n490, n489, n488};
  assign n498 = {n496, n497};
  /* fppowbf16.vhdl:3586:70  */
  assign n499 = {n498, logf_normal};
  /* fppowbf16.vhdl:3588:40  */
  assign n500 = ~sr_d6;
  /* fppowbf16.vhdl:3588:30  */
  assign n501 = n500 ? logf_normal_pad : n502;
  /* fppowbf16.vhdl:3588:50  */
  assign n502 = ~logf_normal_pad;
  /* fppowbf16.vhdl:3589:4  */
  intadder_38_freq500_uid51 lnadder (
    .clk(clk),
    .x(lnaddx),
    .y(lnaddy),
    .cin(sr),
    .r(lnadder_n503));
  /* fppowbf16.vhdl:3595:4  */
  normalizer_z_38_30_16_freq500_uid53 final_norm (
    .clk(clk),
    .x(log_normal),
    .count(final_norm_n506),
    .r(final_norm_n507));
  /* fppowbf16.vhdl:3600:36  */
  assign n512 = z2o2_full_dummy[27:14]; // extract
  /* fppowbf16.vhdl:3601:4  */
  rightshifter14_by_max_13_freq500_uid55 ao_rshift (
    .clk(clk),
    .x(z2o2_small_bs),
    .s(shiftvalinr),
    .r(ao_rshift_n513));
  /* fppowbf16.vhdl:3607:61  */
  assign n516 = z2o2_small_s[26:13]; // extract
  /* fppowbf16.vhdl:3607:47  */
  assign n518 = {9'b000000000, n516};
  /* fppowbf16.vhdl:3609:33  */
  assign n520 = {small_absz0_normd, 13'b0000000000000};
  /* fppowbf16.vhdl:3610:29  */
  assign n521 = sr_d6 ? z2o2_small : n522;
  /* fppowbf16.vhdl:3610:49  */
  assign n522 = ~z2o2_small;
  /* fppowbf16.vhdl:3611:14  */
  assign n523 = ~sr;
  /* fppowbf16.vhdl:3612:4  */
  intadder_23_freq500_uid57 log_small_adder (
    .clk(clk),
    .x(z_small),
    .y(log_smally),
    .cin(nsrcin),
    .r(log_small_adder_n524));
  /* fppowbf16.vhdl:3619:35  */
  assign n528 = log_small[22]; // extract
  /* fppowbf16.vhdl:3619:21  */
  assign n529 = n528 ? 2'b11 : n534;
  /* fppowbf16.vhdl:3620:35  */
  assign n531 = log_small[22:21]; // extract
  /* fppowbf16.vhdl:3620:56  */
  assign n533 = n531 == 2'b01;
  /* fppowbf16.vhdl:3620:11  */
  assign n534 = n533 ? 2'b10 : 2'b01;
  /* fppowbf16.vhdl:3626:46  */
  assign n538 = {6'b011111, e0_sub};
  /* fppowbf16.vhdl:3626:84  */
  assign n540 = {3'b000, lzo_d3};
  /* fppowbf16.vhdl:3626:57  */
  assign n541 = n538 - n540;
  /* fppowbf16.vhdl:3627:32  */
  assign n542 = log_small[22:2]; // extract
  /* fppowbf16.vhdl:3627:64  */
  assign n543 = log_small[22]; // extract
  /* fppowbf16.vhdl:3627:50  */
  assign n544 = n543 ? n542 : n547;
  /* fppowbf16.vhdl:3628:26  */
  assign n545 = log_small[21:1]; // extract
  /* fppowbf16.vhdl:3628:57  */
  assign n546 = log_small[21]; // extract
  /* fppowbf16.vhdl:3628:12  */
  assign n547 = n546 ? n545 : n548;
  /* fppowbf16.vhdl:3629:26  */
  assign n548 = log_small[20:0]; // extract
  /* fppowbf16.vhdl:3631:33  */
  assign n550 = small_d6 ? e_small_d4 : n553;
  /* fppowbf16.vhdl:3632:48  */
  assign n552 = {3'b000, e_normal};
  /* fppowbf16.vhdl:3632:25  */
  assign n553 = e0offset_d10 - n552;
  /* fppowbf16.vhdl:3633:32  */
  assign n554 = log_small_normd_d5[19:0]; // extract
  /* fppowbf16.vhdl:3633:50  */
  assign n556 = {n554, 1'b0};
  /* fppowbf16.vhdl:3633:56  */
  assign n557 = small_d7 ? n556 : n558;
  /* fppowbf16.vhdl:3634:28  */
  assign n558 = log_normal_normd[28:8]; // extract
  /* fppowbf16.vhdl:3635:18  */
  assign n559 = log_g[3]; // extract
  /* fppowbf16.vhdl:3637:26  */
  assign n560 = log_g[20:4]; // extract
  /* fppowbf16.vhdl:3637:19  */
  assign n561 = {er_d1, n560};
  /* fppowbf16.vhdl:3638:39  */
  assign n563 = {24'b000000000000000000000000, round};
  /* fppowbf16.vhdl:3639:4  */
  intadder_25_freq500_uid60 finalroundadder (
    .clk(clk),
    .x(frax),
    .y(fray),
    .cin(n564),
    .r(finalroundadder_n565));
  /* fppowbf16.vhdl:3645:36  */
  assign n569 = xexnsgn_d11[2]; // extract
  /* fppowbf16.vhdl:3645:56  */
  assign n570 = xexnsgn_d11[1]; // extract
  /* fppowbf16.vhdl:3645:74  */
  assign n571 = xexnsgn_d11[0]; // extract
  /* fppowbf16.vhdl:3645:60  */
  assign n572 = n570 | n571;
  /* fppowbf16.vhdl:3645:40  */
  assign n573 = n569 & n572;
  /* fppowbf16.vhdl:3645:95  */
  assign n574 = xexnsgn_d11[1]; // extract
  /* fppowbf16.vhdl:3645:114  */
  assign n575 = xexnsgn_d11[0]; // extract
  /* fppowbf16.vhdl:3645:99  */
  assign n576 = n574 & n575;
  /* fppowbf16.vhdl:3645:80  */
  assign n577 = n573 | n576;
  /* fppowbf16.vhdl:3645:18  */
  assign n578 = n577 ? 3'b110 : n583;
  /* fppowbf16.vhdl:3646:53  */
  assign n580 = xexnsgn_d11[2:1]; // extract
  /* fppowbf16.vhdl:3646:66  */
  assign n582 = n580 == 2'b00;
  /* fppowbf16.vhdl:3645:126  */
  assign n583 = n582 ? 3'b101 : n588;
  /* fppowbf16.vhdl:3647:53  */
  assign n585 = xexnsgn_d11[2:1]; // extract
  /* fppowbf16.vhdl:3647:66  */
  assign n587 = n585 == 2'b10;
  /* fppowbf16.vhdl:3646:74  */
  assign n588 = n587 ? 3'b100 : n601;
  /* fppowbf16.vhdl:3648:36  */
  assign n590 = {2'b00, sr_d11};
  /* fppowbf16.vhdl:3648:69  */
  assign n591 = log_normal_normd[29]; // extract
  /* fppowbf16.vhdl:3648:83  */
  assign n592 = ~n591;
  /* fppowbf16.vhdl:3648:102  */
  assign n593 = ~small_d7;
  /* fppowbf16.vhdl:3648:89  */
  assign n594 = n593 & n592;
  /* fppowbf16.vhdl:3648:134  */
  assign n595 = log_small_normd_d5[20]; // extract
  /* fppowbf16.vhdl:3648:142  */
  assign n596 = ~n595;
  /* fppowbf16.vhdl:3648:148  */
  assign n597 = small_d7 & n596;
  /* fppowbf16.vhdl:3648:109  */
  assign n598 = n594 | n597;
  /* fppowbf16.vhdl:3648:187  */
  assign n599 = small_d7 & ufl_d11;
  /* fppowbf16.vhdl:3648:169  */
  assign n600 = n598 | n599;
  /* fppowbf16.vhdl:3647:74  */
  assign n601 = n600 ? n590 : n603;
  /* fppowbf16.vhdl:3649:37  */
  assign n603 = {2'b01, sr_d11};
  /* fppowbf16.vhdl:3650:14  */
  assign n604 = {rexn, efr};
  /* fppowbf16.vhdl:3398:10  */
  always @(posedge clk)
    n605 <= xexnsgn;
  /* fppowbf16.vhdl:3398:10  */
  always @(posedge clk)
    n606 <= xexnsgn_d1;
  /* fppowbf16.vhdl:3398:10  */
  always @(posedge clk)
    n607 <= xexnsgn_d2;
  /* fppowbf16.vhdl:3398:10  */
  always @(posedge clk)
    n608 <= xexnsgn_d3;
  /* fppowbf16.vhdl:3398:10  */
  always @(posedge clk)
    n609 <= xexnsgn_d4;
  /* fppowbf16.vhdl:3398:10  */
  always @(posedge clk)
    n610 <= xexnsgn_d5;
  /* fppowbf16.vhdl:3398:10  */
  always @(posedge clk)
    n611 <= xexnsgn_d6;
  /* fppowbf16.vhdl:3398:10  */
  always @(posedge clk)
    n612 <= xexnsgn_d7;
  /* fppowbf16.vhdl:3398:10  */
  always @(posedge clk)
    n613 <= xexnsgn_d8;
  /* fppowbf16.vhdl:3398:10  */
  always @(posedge clk)
    n614 <= xexnsgn_d9;
  /* fppowbf16.vhdl:3398:10  */
  always @(posedge clk)
    n615 <= xexnsgn_d10;
  /* fppowbf16.vhdl:3398:10  */
  always @(posedge clk)
    n616 <= y0;
  /* fppowbf16.vhdl:3398:10  */
  always @(posedge clk)
    n617 <= sr;
  /* fppowbf16.vhdl:3398:10  */
  always @(posedge clk)
    n618 <= sr_d1;
  /* fppowbf16.vhdl:3398:10  */
  always @(posedge clk)
    n619 <= sr_d2;
  /* fppowbf16.vhdl:3398:10  */
  always @(posedge clk)
    n620 <= sr_d3;
  /* fppowbf16.vhdl:3398:10  */
  always @(posedge clk)
    n621 <= sr_d4;
  /* fppowbf16.vhdl:3398:10  */
  always @(posedge clk)
    n622 <= sr_d5;
  /* fppowbf16.vhdl:3398:10  */
  always @(posedge clk)
    n623 <= sr_d6;
  /* fppowbf16.vhdl:3398:10  */
  always @(posedge clk)
    n624 <= sr_d7;
  /* fppowbf16.vhdl:3398:10  */
  always @(posedge clk)
    n625 <= sr_d8;
  /* fppowbf16.vhdl:3398:10  */
  always @(posedge clk)
    n626 <= sr_d9;
  /* fppowbf16.vhdl:3398:10  */
  always @(posedge clk)
    n627 <= sr_d10;
  /* fppowbf16.vhdl:3398:10  */
  always @(posedge clk)
    n628 <= eeqzero;
  /* fppowbf16.vhdl:3398:10  */
  always @(posedge clk)
    n629 <= eeqzero_d1;
  /* fppowbf16.vhdl:3398:10  */
  always @(posedge clk)
    n630 <= eeqzero_d2;
  /* fppowbf16.vhdl:3398:10  */
  always @(posedge clk)
    n631 <= eeqzero_d3;
  /* fppowbf16.vhdl:3398:10  */
  always @(posedge clk)
    n632 <= lzo;
  /* fppowbf16.vhdl:3398:10  */
  always @(posedge clk)
    n633 <= lzo_d1;
  /* fppowbf16.vhdl:3398:10  */
  always @(posedge clk)
    n634 <= lzo_d2;
  /* fppowbf16.vhdl:3398:10  */
  always @(posedge clk)
    n635 <= pfinal_s;
  /* fppowbf16.vhdl:3398:10  */
  always @(posedge clk)
    n636 <= pfinal_s_d1;
  /* fppowbf16.vhdl:3398:10  */
  always @(posedge clk)
    n637 <= pfinal_s_d2;
  /* fppowbf16.vhdl:3398:10  */
  always @(posedge clk)
    n638 <= dorr;
  /* fppowbf16.vhdl:3398:10  */
  always @(posedge clk)
    n639 <= dorr_d1;
  /* fppowbf16.vhdl:3398:10  */
  always @(posedge clk)
    n640 <= \small ;
  /* fppowbf16.vhdl:3398:10  */
  always @(posedge clk)
    n641 <= small_d1;
  /* fppowbf16.vhdl:3398:10  */
  always @(posedge clk)
    n642 <= small_d2;
  /* fppowbf16.vhdl:3398:10  */
  always @(posedge clk)
    n643 <= small_d3;
  /* fppowbf16.vhdl:3398:10  */
  always @(posedge clk)
    n644 <= small_d4;
  /* fppowbf16.vhdl:3398:10  */
  always @(posedge clk)
    n645 <= small_d5;
  /* fppowbf16.vhdl:3398:10  */
  always @(posedge clk)
    n646 <= small_d6;
  /* fppowbf16.vhdl:3398:10  */
  always @(posedge clk)
    n647 <= small_absz0_normd;
  /* fppowbf16.vhdl:3398:10  */
  always @(posedge clk)
    n648 <= inva0;
  /* fppowbf16.vhdl:3398:10  */
  always @(posedge clk)
    n649 <= a1;
  /* fppowbf16.vhdl:3398:10  */
  always @(posedge clk)
    n650 <= zm1;
  /* fppowbf16.vhdl:3398:10  */
  always @(posedge clk)
    n651 <= zfinal;
  /* fppowbf16.vhdl:3398:10  */
  always @(posedge clk)
    n652 <= zfinal_d1;
  /* fppowbf16.vhdl:3398:10  */
  always @(posedge clk)
    n653 <= ufl;
  /* fppowbf16.vhdl:3398:10  */
  always @(posedge clk)
    n654 <= ufl_d1;
  /* fppowbf16.vhdl:3398:10  */
  always @(posedge clk)
    n655 <= ufl_d2;
  /* fppowbf16.vhdl:3398:10  */
  always @(posedge clk)
    n656 <= ufl_d3;
  /* fppowbf16.vhdl:3398:10  */
  always @(posedge clk)
    n657 <= ufl_d4;
  /* fppowbf16.vhdl:3398:10  */
  always @(posedge clk)
    n658 <= ufl_d5;
  /* fppowbf16.vhdl:3398:10  */
  always @(posedge clk)
    n659 <= ufl_d6;
  /* fppowbf16.vhdl:3398:10  */
  always @(posedge clk)
    n660 <= ufl_d7;
  /* fppowbf16.vhdl:3398:10  */
  always @(posedge clk)
    n661 <= ufl_d8;
  /* fppowbf16.vhdl:3398:10  */
  always @(posedge clk)
    n662 <= ufl_d9;
  /* fppowbf16.vhdl:3398:10  */
  always @(posedge clk)
    n663 <= ufl_d10;
  /* fppowbf16.vhdl:3398:10  */
  always @(posedge clk)
    n664 <= e_small;
  /* fppowbf16.vhdl:3398:10  */
  always @(posedge clk)
    n665 <= e_small_d1;
  /* fppowbf16.vhdl:3398:10  */
  always @(posedge clk)
    n666 <= e_small_d2;
  /* fppowbf16.vhdl:3398:10  */
  always @(posedge clk)
    n667 <= e_small_d3;
  /* fppowbf16.vhdl:3398:10  */
  always @(posedge clk)
    n668 <= log_small_normd;
  /* fppowbf16.vhdl:3398:10  */
  always @(posedge clk)
    n669 <= log_small_normd_d1;
  /* fppowbf16.vhdl:3398:10  */
  always @(posedge clk)
    n670 <= log_small_normd_d2;
  /* fppowbf16.vhdl:3398:10  */
  always @(posedge clk)
    n671 <= log_small_normd_d3;
  /* fppowbf16.vhdl:3398:10  */
  always @(posedge clk)
    n672 <= log_small_normd_d4;
  /* fppowbf16.vhdl:3398:10  */
  always @(posedge clk)
    n673 <= e0offset;
  /* fppowbf16.vhdl:3398:10  */
  always @(posedge clk)
    n674 <= e0offset_d1;
  /* fppowbf16.vhdl:3398:10  */
  always @(posedge clk)
    n675 <= e0offset_d2;
  /* fppowbf16.vhdl:3398:10  */
  always @(posedge clk)
    n676 <= e0offset_d3;
  /* fppowbf16.vhdl:3398:10  */
  always @(posedge clk)
    n677 <= e0offset_d4;
  /* fppowbf16.vhdl:3398:10  */
  always @(posedge clk)
    n678 <= e0offset_d5;
  /* fppowbf16.vhdl:3398:10  */
  always @(posedge clk)
    n679 <= e0offset_d6;
  /* fppowbf16.vhdl:3398:10  */
  always @(posedge clk)
    n680 <= e0offset_d7;
  /* fppowbf16.vhdl:3398:10  */
  always @(posedge clk)
    n681 <= e0offset_d8;
  /* fppowbf16.vhdl:3398:10  */
  always @(posedge clk)
    n682 <= e0offset_d9;
  /* fppowbf16.vhdl:3398:10  */
  always @(posedge clk)
    n683 <= er;
endmodule

module lzc_7_freq500_uid7
  (input  clk,
   input  [6:0] i,
   output [2:0] o);
  wire [6:0] level3;
  wire digit2;
  wire [2:0] level2;
  wire [1:0] lowbits;
  wire outhighbits;
  wire [3:0] n247;
  wire n249;
  wire n250;
  wire [2:0] n252;
  wire [2:0] n253;
  wire [2:0] n254;
  wire n257;
  wire n260;
  wire n263;
  wire n266;
  wire [3:0] n268;
  reg [1:0] n269;
  wire [2:0] n271;
  assign o = n271; //(module output)
  /* fppowbf16.vhdl:1951:26  */
  assign digit2 = n250; // (signal)
  /* fppowbf16.vhdl:1932:8  */
  assign level2 = n253; // (signal)
  /* fppowbf16.vhdl:1934:8  */
  assign lowbits = n269; // (signal)
  /* fppowbf16.vhdl:1936:8  */
  assign outhighbits = digit2; // (signal)
  /* fppowbf16.vhdl:1942:28  */
  assign n247 = level3[6:3]; // extract
  /* fppowbf16.vhdl:1942:41  */
  assign n249 = n247 == 4'b0000;
  /* fppowbf16.vhdl:1942:17  */
  assign n250 = n249 ? 1'b1 : 1'b0;
  /* fppowbf16.vhdl:1943:19  */
  assign n252 = level3[2:0]; // extract
  /* fppowbf16.vhdl:1943:32  */
  assign n253 = digit2 ? n252 : n254;
  /* fppowbf16.vhdl:1943:59  */
  assign n254 = level3[6:4]; // extract
  /* fppowbf16.vhdl:1946:12  */
  assign n257 = level2 == 3'b000;
  /* fppowbf16.vhdl:1947:12  */
  assign n260 = level2 == 3'b001;
  /* fppowbf16.vhdl:1948:12  */
  assign n263 = level2 == 3'b010;
  /* fppowbf16.vhdl:1949:12  */
  assign n266 = level2 == 3'b011;
  assign n268 = {n266, n263, n260, n257};
  /* fppowbf16.vhdl:1945:4  */
  always @*
    case (n268)
      4'b1000: n269 = 2'b01;
      4'b0100: n269 = 2'b01;
      4'b0010: n269 = 2'b10;
      4'b0001: n269 = 2'b11;
      default: n269 = 2'b00;
    endcase
  /* fppowbf16.vhdl:1952:21  */
  assign n271 = {outhighbits, lowbits};
endmodule

module intadder_16_freq500_uid5
  (input  clk,
   input  [15:0] x,
   input  [15:0] y,
   input  cin,
   output [15:0] r);
  wire [15:0] rtmp;
  wire [15:0] n242;
  wire [15:0] n243;
  wire [15:0] n244;
  assign r = rtmp; //(module output)
  /* fppowbf16.vhdl:1891:8  */
  assign rtmp = n244; // (signal)
  /* fppowbf16.vhdl:1894:14  */
  assign n242 = x + y;
  /* fppowbf16.vhdl:1894:18  */
  assign n243 = {15'b0, cin};  //  uext
  /* fppowbf16.vhdl:1894:18  */
  assign n244 = n242 + n243;
endmodule

module top_module
  (input  clk,
   input  [17:0] X,
   input  [17:0] Y,
   output [17:0] R);
  wire [1:0] flagsx;
  wire signx;
  wire signx_d1;
  wire [7:0] expfieldx;
  wire [6:0] fracx;
  wire [1:0] flagsy;
  wire signy;
  wire signy_d1;
  wire signy_d2;
  wire [7:0] expfieldy;
  wire [6:0] fracy;
  wire zerox;
  wire zerox_d1;
  wire zerox_d2;
  wire zeroy;
  wire zeroy_d1;
  wire normalx;
  wire normalx_d1;
  wire normaly;
  wire normaly_d1;
  wire normaly_d2;
  wire infx;
  wire infx_d1;
  wire infx_d2;
  wire infy;
  wire infy_d1;
  wire infy_d2;
  wire s_nan_in;
  wire s_nan_in_d1;
  wire [14:0] oneexpfrac;
  wire [15:0] expfracx;
  wire [15:0] oneexpfraccompl;
  wire [15:0] cmpxoneres;
  wire xisoneandnormal;
  wire absxgtoneandnormal;
  wire absxgtoneandnormal_d1;
  wire absxgtoneandnormal_d2;
  wire absxltoneandnormal;
  wire absxltoneandnormal_d1;
  wire absxltoneandnormal_d2;
  wire [6:0] fracyreverted;
  wire [2:0] z_righty;
  wire [2:0] z_righty_d1;
  wire [8:0] weightlsbypre;
  wire [8:0] weightlsbypre_d1;
  wire [8:0] weightlsby;
  wire [8:0] weightlsby_d1;
  wire oddinty;
  wire oddinty_d1;
  wire eveninty;
  wire notintnormaly;
  wire risinfspecialcase;
  wire riszerospecialcase;
  wire risone;
  wire risnan;
  wire signr;
  wire [27:0] login;
  wire [27:0] lnx;
  wire [28:0] p;
  wire [17:0] e;
  wire [1:0] flagse;
  wire riszerofromexp;
  wire riszero;
  wire risinffromexp;
  wire risinf;
  wire [1:0] flagr;
  wire [14:0] r_expfrac;
  wire [1:0] n27;
  wire n28;
  wire [7:0] n29;
  wire [6:0] n30;
  wire [1:0] n31;
  wire n32;
  wire [7:0] n33;
  wire [6:0] n34;
  wire n37;
  wire n38;
  wire n42;
  wire n43;
  wire n47;
  wire n48;
  wire n52;
  wire n53;
  wire n57;
  wire n58;
  wire n62;
  wire n63;
  wire n67;
  wire n69;
  wire n70;
  wire n71;
  wire [8:0] n75;
  wire [15:0] n76;
  wire [14:0] n77;
  wire [15:0] n79;
  localparam n80 = 1'b1;
  wire [15:0] cmpxone_n81;
  wire [17:0] n86;
  wire n87;
  wire n88;
  wire n90;
  wire n91;
  wire n92;
  wire n93;
  wire n94;
  wire n95;
  wire n96;
  wire n97;
  wire n98;
  wire [1:0] n99;
  wire n100;
  wire [2:0] n101;
  wire n102;
  wire [3:0] n103;
  wire n104;
  wire [4:0] n105;
  wire n106;
  wire [5:0] n107;
  wire n108;
  wire [6:0] n109;
  wire [2:0] fppow_8_7_freq500_uid2right1counter_n110;
  wire [8:0] n114;
  wire [8:0] n116;
  wire [8:0] n117;
  wire [8:0] n118;
  wire n120;
  wire n121;
  wire n123;
  wire n124;
  wire n125;
  wire n126;
  wire n127;
  wire n129;
  wire n130;
  wire n132;
  wire n133;
  wire n134;
  wire n135;
  wire n136;
  wire n137;
  wire n138;
  wire n139;
  wire n140;
  wire n141;
  wire n142;
  wire n143;
  wire n144;
  wire n145;
  wire n146;
  wire n147;
  wire n148;
  wire n149;
  wire n150;
  wire n151;
  wire n152;
  wire n153;
  wire n154;
  wire n155;
  wire n156;
  wire n157;
  wire n158;
  wire n159;
  wire n160;
  wire n161;
  wire n162;
  wire n163;
  wire n164;
  wire n165;
  wire n166;
  wire n167;
  wire n168;
  wire n169;
  wire n170;
  wire n171;
  wire n172;
  wire n173;
  wire n174;
  wire n175;
  wire n176;
  wire n177;
  wire n178;
  wire [2:0] n180;
  wire [10:0] n181;
  wire [17:0] n182;
  wire [27:0] n184;
  wire [27:0] fppow_8_7_freq500_uid2log_n185;
  wire [28:0] fppow_8_7_freq500_uid2mult_n188;
  wire [17:0] fppow_8_7_freq500_uid2exp_n191;
  wire [1:0] n194;
  wire n197;
  wire n198;
  wire n200;
  wire n203;
  wire n204;
  wire n206;
  wire [1:0] n208;
  wire [1:0] n210;
  wire [1:0] n212;
  wire [14:0] n215;
  wire [14:0] n216;
  wire [2:0] n217;
  wire [17:0] n218;
  reg n219;
  reg n220;
  reg n221;
  reg n222;
  reg n223;
  reg n224;
  reg n225;
  reg n226;
  reg n227;
  reg n228;
  reg n229;
  reg n230;
  reg n231;
  reg n232;
  reg n233;
  reg n234;
  reg n235;
  reg n236;
  reg [2:0] n237;
  reg [8:0] n238;
  reg [8:0] n239;
  reg n240;
  assign R = n218; //(module output)
  /* fppowbf16.vhdl:5031:8  */
  assign flagsx = n27; // (signal)
  /* fppowbf16.vhdl:5033:8  */
  assign signx = n28; // (signal)
  /* fppowbf16.vhdl:5033:15  */
  assign signx_d1 = n219; // (signal)
  /* fppowbf16.vhdl:5035:8  */
  assign expfieldx = n29; // (signal)
  /* fppowbf16.vhdl:5037:8  */
  assign fracx = n30; // (signal)
  /* fppowbf16.vhdl:5039:8  */
  assign flagsy = n31; // (signal)
  /* fppowbf16.vhdl:5041:8  */
  assign signy = n32; // (signal)
  /* fppowbf16.vhdl:5041:15  */
  assign signy_d1 = n220; // (signal)
  /* fppowbf16.vhdl:5041:25  */
  assign signy_d2 = n221; // (signal)
  /* fppowbf16.vhdl:5043:8  */
  assign expfieldy = n33; // (signal)
  /* fppowbf16.vhdl:5045:8  */
  assign fracy = n34; // (signal)
  /* fppowbf16.vhdl:5047:8  */
  assign zerox = n38; // (signal)
  /* fppowbf16.vhdl:5047:15  */
  assign zerox_d1 = n222; // (signal)
  /* fppowbf16.vhdl:5047:25  */
  assign zerox_d2 = n223; // (signal)
  /* fppowbf16.vhdl:5049:8  */
  assign zeroy = n43; // (signal)
  /* fppowbf16.vhdl:5049:15  */
  assign zeroy_d1 = n224; // (signal)
  /* fppowbf16.vhdl:5051:8  */
  assign normalx = n48; // (signal)
  /* fppowbf16.vhdl:5051:17  */
  assign normalx_d1 = n225; // (signal)
  /* fppowbf16.vhdl:5053:8  */
  assign normaly = n53; // (signal)
  /* fppowbf16.vhdl:5053:17  */
  assign normaly_d1 = n226; // (signal)
  /* fppowbf16.vhdl:5053:29  */
  assign normaly_d2 = n227; // (signal)
  /* fppowbf16.vhdl:5055:8  */
  assign infx = n58; // (signal)
  /* fppowbf16.vhdl:5055:14  */
  assign infx_d1 = n228; // (signal)
  /* fppowbf16.vhdl:5055:23  */
  assign infx_d2 = n229; // (signal)
  /* fppowbf16.vhdl:5057:8  */
  assign infy = n63; // (signal)
  /* fppowbf16.vhdl:5057:14  */
  assign infy_d1 = n230; // (signal)
  /* fppowbf16.vhdl:5057:23  */
  assign infy_d2 = n231; // (signal)
  /* fppowbf16.vhdl:5059:8  */
  assign s_nan_in = n71; // (signal)
  /* fppowbf16.vhdl:5059:18  */
  assign s_nan_in_d1 = n232; // (signal)
  /* fppowbf16.vhdl:5061:8  */
  assign oneexpfrac = 15'b011111110000000; // (signal)
  /* fppowbf16.vhdl:5063:8  */
  assign expfracx = n76; // (signal)
  /* fppowbf16.vhdl:5065:8  */
  assign oneexpfraccompl = n79; // (signal)
  /* fppowbf16.vhdl:5067:8  */
  assign cmpxoneres = cmpxone_n81; // (signal)
  /* fppowbf16.vhdl:5069:8  */
  assign xisoneandnormal = n88; // (signal)
  /* fppowbf16.vhdl:5071:8  */
  assign absxgtoneandnormal = n94; // (signal)
  /* fppowbf16.vhdl:5071:28  */
  assign absxgtoneandnormal_d1 = n233; // (signal)
  /* fppowbf16.vhdl:5071:51  */
  assign absxgtoneandnormal_d2 = n234; // (signal)
  /* fppowbf16.vhdl:5073:8  */
  assign absxltoneandnormal = n96; // (signal)
  /* fppowbf16.vhdl:5073:28  */
  assign absxltoneandnormal_d1 = n235; // (signal)
  /* fppowbf16.vhdl:5073:51  */
  assign absxltoneandnormal_d2 = n236; // (signal)
  /* fppowbf16.vhdl:5075:8  */
  assign fracyreverted = n109; // (signal)
  /* fppowbf16.vhdl:5077:8  */
  assign z_righty = fppow_8_7_freq500_uid2right1counter_n110; // (signal)
  /* fppowbf16.vhdl:5077:18  */
  assign z_righty_d1 = n237; // (signal)
  /* fppowbf16.vhdl:5079:8  */
  assign weightlsbypre = n116; // (signal)
  /* fppowbf16.vhdl:5079:23  */
  assign weightlsbypre_d1 = n238; // (signal)
  /* fppowbf16.vhdl:5081:8  */
  assign weightlsby = n118; // (signal)
  /* fppowbf16.vhdl:5081:20  */
  assign weightlsby_d1 = n239; // (signal)
  /* fppowbf16.vhdl:5083:8  */
  assign oddinty = n121; // (signal)
  /* fppowbf16.vhdl:5083:17  */
  assign oddinty_d1 = n240; // (signal)
  /* fppowbf16.vhdl:5085:8  */
  assign eveninty = n127; // (signal)
  /* fppowbf16.vhdl:5087:8  */
  assign notintnormaly = n130; // (signal)
  /* fppowbf16.vhdl:5089:8  */
  assign risinfspecialcase = n148; // (signal)
  /* fppowbf16.vhdl:5091:8  */
  assign riszerospecialcase = n166; // (signal)
  /* fppowbf16.vhdl:5093:8  */
  assign risone = n172; // (signal)
  /* fppowbf16.vhdl:5095:8  */
  assign risnan = n177; // (signal)
  /* fppowbf16.vhdl:5097:8  */
  assign signr = n178; // (signal)
  /* fppowbf16.vhdl:5099:8  */
  assign login = n184; // (signal)
  /* fppowbf16.vhdl:5101:8  */
  assign lnx = fppow_8_7_freq500_uid2log_n185; // (signal)
  /* fppowbf16.vhdl:5103:8  */
  assign p = fppow_8_7_freq500_uid2mult_n188; // (signal)
  /* fppowbf16.vhdl:5105:8  */
  assign e = fppow_8_7_freq500_uid2exp_n191; // (signal)
  /* fppowbf16.vhdl:5107:8  */
  assign flagse = n194; // (signal)
  /* fppowbf16.vhdl:5109:8  */
  assign riszerofromexp = n198; // (signal)
  /* fppowbf16.vhdl:5111:8  */
  assign riszero = n200; // (signal)
  /* fppowbf16.vhdl:5113:8  */
  assign risinffromexp = n204; // (signal)
  /* fppowbf16.vhdl:5115:8  */
  assign risinf = n206; // (signal)
  /* fppowbf16.vhdl:5117:8  */
  assign flagr = n208; // (signal)
  /* fppowbf16.vhdl:5119:8  */
  assign r_expfrac = n215; // (signal)
  /* fppowbf16.vhdl:5151:15  */
  assign n27 = X[17:16]; // extract
  /* fppowbf16.vhdl:5152:14  */
  assign n28 = X[15]; // extract
  /* fppowbf16.vhdl:5153:18  */
  assign n29 = X[14:7]; // extract
  /* fppowbf16.vhdl:5154:14  */
  assign n30 = X[6:0]; // extract
  /* fppowbf16.vhdl:5155:15  */
  assign n31 = Y[17:16]; // extract
  /* fppowbf16.vhdl:5156:14  */
  assign n32 = Y[15]; // extract
  /* fppowbf16.vhdl:5157:18  */
  assign n33 = Y[14:7]; // extract
  /* fppowbf16.vhdl:5158:14  */
  assign n34 = Y[6:0]; // extract
  /* fppowbf16.vhdl:5161:28  */
  assign n37 = flagsx == 2'b00;
  /* fppowbf16.vhdl:5161:17  */
  assign n38 = n37 ? 1'b1 : 1'b0;
  /* fppowbf16.vhdl:5162:28  */
  assign n42 = flagsy == 2'b00;
  /* fppowbf16.vhdl:5162:17  */
  assign n43 = n42 ? 1'b1 : 1'b0;
  /* fppowbf16.vhdl:5164:30  */
  assign n47 = flagsx == 2'b01;
  /* fppowbf16.vhdl:5164:19  */
  assign n48 = n47 ? 1'b1 : 1'b0;
  /* fppowbf16.vhdl:5165:30  */
  assign n52 = flagsy == 2'b01;
  /* fppowbf16.vhdl:5165:19  */
  assign n53 = n52 ? 1'b1 : 1'b0;
  /* fppowbf16.vhdl:5167:27  */
  assign n57 = flagsx == 2'b10;
  /* fppowbf16.vhdl:5167:16  */
  assign n58 = n57 ? 1'b1 : 1'b0;
  /* fppowbf16.vhdl:5168:27  */
  assign n62 = flagsy == 2'b10;
  /* fppowbf16.vhdl:5168:16  */
  assign n63 = n62 ? 1'b1 : 1'b0;
  /* fppowbf16.vhdl:5170:31  */
  assign n67 = flagsx == 2'b11;
  /* fppowbf16.vhdl:5170:46  */
  assign n69 = flagsy == 2'b11;
  /* fppowbf16.vhdl:5170:37  */
  assign n70 = n67 | n69;
  /* fppowbf16.vhdl:5170:20  */
  assign n71 = n70 ? 1'b1 : 1'b0;
  /* fppowbf16.vhdl:5173:19  */
  assign n75 = {1'b0, expfieldx};
  /* fppowbf16.vhdl:5173:31  */
  assign n76 = {n75, fracx};
  /* fppowbf16.vhdl:5174:30  */
  assign n77 = ~oneexpfrac;
  /* fppowbf16.vhdl:5174:27  */
  assign n79 = {1'b1, n77};
  /* fppowbf16.vhdl:5175:4  */
  intadder_16_freq500_uid5 cmpxone (
    .clk(clk),
    .x(expfracx),
    .y(oneexpfraccompl),
    .cin(n80),
    .r(cmpxone_n81));
  /* fppowbf16.vhdl:5181:43  */
  assign n86 = {3'b010, oneexpfrac};
  /* fppowbf16.vhdl:5181:34  */
  assign n87 = X == n86;
  /* fppowbf16.vhdl:5181:27  */
  assign n88 = n87 ? 1'b1 : 1'b0;
  /* fppowbf16.vhdl:5182:39  */
  assign n90 = ~xisoneandnormal;
  /* fppowbf16.vhdl:5182:34  */
  assign n91 = normalx & n90;
  /* fppowbf16.vhdl:5182:79  */
  assign n92 = cmpxoneres[15]; // extract
  /* fppowbf16.vhdl:5182:65  */
  assign n93 = ~n92;
  /* fppowbf16.vhdl:5182:60  */
  assign n94 = n91 & n93;
  /* fppowbf16.vhdl:5183:48  */
  assign n95 = cmpxoneres[15]; // extract
  /* fppowbf16.vhdl:5183:34  */
  assign n96 = normalx & n95;
  /* fppowbf16.vhdl:5184:26  */
  assign n97 = fracy[0]; // extract
  /* fppowbf16.vhdl:5184:35  */
  assign n98 = fracy[1]; // extract
  /* fppowbf16.vhdl:5184:29  */
  assign n99 = {n97, n98};
  /* fppowbf16.vhdl:5184:44  */
  assign n100 = fracy[2]; // extract
  /* fppowbf16.vhdl:5184:38  */
  assign n101 = {n99, n100};
  /* fppowbf16.vhdl:5184:53  */
  assign n102 = fracy[3]; // extract
  /* fppowbf16.vhdl:5184:47  */
  assign n103 = {n101, n102};
  /* fppowbf16.vhdl:5184:62  */
  assign n104 = fracy[4]; // extract
  /* fppowbf16.vhdl:5184:56  */
  assign n105 = {n103, n104};
  /* fppowbf16.vhdl:5184:71  */
  assign n106 = fracy[5]; // extract
  /* fppowbf16.vhdl:5184:65  */
  assign n107 = {n105, n106};
  /* fppowbf16.vhdl:5184:80  */
  assign n108 = fracy[6]; // extract
  /* fppowbf16.vhdl:5184:74  */
  assign n109 = {n107, n108};
  /* fppowbf16.vhdl:5185:4  */
  lzc_7_freq500_uid7 fppow_8_7_freq500_uid2right1counter (
    .clk(clk),
    .i(fracyreverted),
    .o(fppow_8_7_freq500_uid2right1counter_n110));
  /* fppowbf16.vhdl:5190:26  */
  assign n114 = {1'b0, expfieldy};
  /* fppowbf16.vhdl:5190:38  */
  assign n116 = n114 - 9'b010000110;
  /* fppowbf16.vhdl:5191:35  */
  assign n117 = {6'b0, z_righty_d1};  //  uext
  /* fppowbf16.vhdl:5191:35  */
  assign n118 = weightlsbypre_d1 + n117;
  /* fppowbf16.vhdl:5192:42  */
  assign n120 = weightlsby == 9'b000000000;
  /* fppowbf16.vhdl:5192:26  */
  assign n121 = n120 ? normaly_d1 : 1'b0;
  /* fppowbf16.vhdl:5193:45  */
  assign n123 = weightlsby_d1[8]; // extract
  /* fppowbf16.vhdl:5193:49  */
  assign n124 = ~n123;
  /* fppowbf16.vhdl:5193:68  */
  assign n125 = ~oddinty_d1;
  /* fppowbf16.vhdl:5193:54  */
  assign n126 = n125 & n124;
  /* fppowbf16.vhdl:5193:27  */
  assign n127 = n126 ? normaly_d2 : 1'b0;
  /* fppowbf16.vhdl:5194:47  */
  assign n129 = weightlsby[8]; // extract
  /* fppowbf16.vhdl:5194:32  */
  assign n130 = n129 ? normaly_d1 : 1'b0;
  /* fppowbf16.vhdl:5198:38  */
  assign n132 = oddinty_d1 | eveninty;
  /* fppowbf16.vhdl:5198:21  */
  assign n133 = zerox_d2 & n132;
  /* fppowbf16.vhdl:5198:52  */
  assign n134 = n133 & signy_d2;
  /* fppowbf16.vhdl:5199:20  */
  assign n135 = zerox_d2 & infy_d2;
  /* fppowbf16.vhdl:5199:32  */
  assign n136 = n135 & signy_d2;
  /* fppowbf16.vhdl:5199:7  */
  assign n137 = n134 | n136;
  /* fppowbf16.vhdl:5200:35  */
  assign n138 = absxgtoneandnormal_d2 & infy_d2;
  /* fppowbf16.vhdl:5200:53  */
  assign n139 = ~signy_d2;
  /* fppowbf16.vhdl:5200:49  */
  assign n140 = n138 & n139;
  /* fppowbf16.vhdl:5200:7  */
  assign n141 = n137 | n140;
  /* fppowbf16.vhdl:5201:35  */
  assign n142 = absxltoneandnormal_d2 & infy_d2;
  /* fppowbf16.vhdl:5201:49  */
  assign n143 = n142 & signy_d2;
  /* fppowbf16.vhdl:5201:7  */
  assign n144 = n141 | n143;
  /* fppowbf16.vhdl:5202:19  */
  assign n145 = infx_d2 & normaly_d2;
  /* fppowbf16.vhdl:5202:40  */
  assign n146 = ~signy_d2;
  /* fppowbf16.vhdl:5202:36  */
  assign n147 = n145 & n146;
  /* fppowbf16.vhdl:5202:7  */
  assign n148 = n144 | n147;
  /* fppowbf16.vhdl:5204:37  */
  assign n149 = oddinty_d1 | eveninty;
  /* fppowbf16.vhdl:5204:20  */
  assign n150 = zerox_d2 & n149;
  /* fppowbf16.vhdl:5204:55  */
  assign n151 = ~signy_d2;
  /* fppowbf16.vhdl:5204:51  */
  assign n152 = n150 & n151;
  /* fppowbf16.vhdl:5205:20  */
  assign n153 = zerox_d2 & infy_d2;
  /* fppowbf16.vhdl:5205:38  */
  assign n154 = ~signy_d2;
  /* fppowbf16.vhdl:5205:34  */
  assign n155 = n153 & n154;
  /* fppowbf16.vhdl:5205:7  */
  assign n156 = n152 | n155;
  /* fppowbf16.vhdl:5206:35  */
  assign n157 = absxltoneandnormal_d2 & infy_d2;
  /* fppowbf16.vhdl:5206:53  */
  assign n158 = ~signy_d2;
  /* fppowbf16.vhdl:5206:49  */
  assign n159 = n157 & n158;
  /* fppowbf16.vhdl:5206:7  */
  assign n160 = n156 | n159;
  /* fppowbf16.vhdl:5207:35  */
  assign n161 = absxgtoneandnormal_d2 & infy_d2;
  /* fppowbf16.vhdl:5207:49  */
  assign n162 = n161 & signy_d2;
  /* fppowbf16.vhdl:5207:7  */
  assign n163 = n160 | n162;
  /* fppowbf16.vhdl:5208:19  */
  assign n164 = infx_d2 & normaly_d2;
  /* fppowbf16.vhdl:5208:36  */
  assign n165 = n164 & signy_d2;
  /* fppowbf16.vhdl:5208:7  */
  assign n166 = n163 | n165;
  /* fppowbf16.vhdl:5211:27  */
  assign n167 = xisoneandnormal & signx;
  /* fppowbf16.vhdl:5211:37  */
  assign n168 = n167 & infy;
  /* fppowbf16.vhdl:5211:7  */
  assign n169 = zeroy | n168;
  /* fppowbf16.vhdl:5212:32  */
  assign n170 = ~signx;
  /* fppowbf16.vhdl:5212:28  */
  assign n171 = xisoneandnormal & n170;
  /* fppowbf16.vhdl:5212:7  */
  assign n172 = n169 | n171;
  /* fppowbf16.vhdl:5213:31  */
  assign n173 = ~zeroy_d1;
  /* fppowbf16.vhdl:5213:27  */
  assign n174 = s_nan_in_d1 & n173;
  /* fppowbf16.vhdl:5213:60  */
  assign n175 = normalx_d1 & signx_d1;
  /* fppowbf16.vhdl:5213:73  */
  assign n176 = n175 & notintnormaly;
  /* fppowbf16.vhdl:5213:45  */
  assign n177 = n174 | n176;
  /* fppowbf16.vhdl:5214:22  */
  assign n178 = signx_d1 & oddinty;
  /* fppowbf16.vhdl:5215:20  */
  assign n180 = {flagsx, 1'b0};
  /* fppowbf16.vhdl:5215:26  */
  assign n181 = {n180, expfieldx};
  /* fppowbf16.vhdl:5215:38  */
  assign n182 = {n181, fracx};
  /* fppowbf16.vhdl:5215:46  */
  assign n184 = {n182, 10'b0000000000};
  /* fppowbf16.vhdl:5216:4  */
  fplogiterative_8_17_0_500_freq500_uid9 fppow_8_7_freq500_uid2log (
    .clk(clk),
    .x(login),
    .r(fppow_8_7_freq500_uid2log_n185));
  /* fppowbf16.vhdl:5220:4  */
  fpmult_8_17_uid62_freq500_uid63 fppow_8_7_freq500_uid2mult (
    .clk(clk),
    .x(lnx),
    .y(Y),
    .r(fppow_8_7_freq500_uid2mult_n188));
  /* fppowbf16.vhdl:5225:4  */
  fpexp_8_7_freq500_uid71 fppow_8_7_freq500_uid2exp (
    .clk(clk),
    .x(p),
    .r(fppow_8_7_freq500_uid2exp_n191));
  /* fppowbf16.vhdl:5229:15  */
  assign n194 = e[17:16]; // extract
  /* fppowbf16.vhdl:5230:37  */
  assign n197 = flagse == 2'b00;
  /* fppowbf16.vhdl:5230:26  */
  assign n198 = n197 ? 1'b1 : 1'b0;
  /* fppowbf16.vhdl:5231:34  */
  assign n200 = riszerospecialcase | riszerofromexp;
  /* fppowbf16.vhdl:5232:37  */
  assign n203 = flagse == 2'b10;
  /* fppowbf16.vhdl:5232:26  */
  assign n204 = n203 ? 1'b1 : 1'b0;
  /* fppowbf16.vhdl:5233:33  */
  assign n206 = risinfspecialcase | risinffromexp;
  /* fppowbf16.vhdl:5235:17  */
  assign n208 = risnan ? 2'b11 : n210;
  /* fppowbf16.vhdl:5236:7  */
  assign n210 = riszero ? 2'b00 : n212;
  /* fppowbf16.vhdl:5237:7  */
  assign n212 = risinf ? 2'b10 : 2'b01;
  /* fppowbf16.vhdl:5239:77  */
  assign n215 = risone ? 15'b011111110000000 : n216;
  /* fppowbf16.vhdl:5240:14  */
  assign n216 = e[14:0]; // extract
  /* fppowbf16.vhdl:5241:15  */
  assign n217 = {flagr, signr};
  /* fppowbf16.vhdl:5241:23  */
  assign n218 = {n217, r_expfrac};
  /* fppowbf16.vhdl:5126:10  */
  always @(posedge clk)
    n219 <= signx;
  /* fppowbf16.vhdl:5126:10  */
  always @(posedge clk)
    n220 <= signy;
  /* fppowbf16.vhdl:5126:10  */
  always @(posedge clk)
    n221 <= signy_d1;
  /* fppowbf16.vhdl:5126:10  */
  always @(posedge clk)
    n222 <= zerox;
  /* fppowbf16.vhdl:5126:10  */
  always @(posedge clk)
    n223 <= zerox_d1;
  /* fppowbf16.vhdl:5126:10  */
  always @(posedge clk)
    n224 <= zeroy;
  /* fppowbf16.vhdl:5126:10  */
  always @(posedge clk)
    n225 <= normalx;
  /* fppowbf16.vhdl:5126:10  */
  always @(posedge clk)
    n226 <= normaly;
  /* fppowbf16.vhdl:5126:10  */
  always @(posedge clk)
    n227 <= normaly_d1;
  /* fppowbf16.vhdl:5126:10  */
  always @(posedge clk)
    n228 <= infx;
  /* fppowbf16.vhdl:5126:10  */
  always @(posedge clk)
    n229 <= infx_d1;
  /* fppowbf16.vhdl:5126:10  */
  always @(posedge clk)
    n230 <= infy;
  /* fppowbf16.vhdl:5126:10  */
  always @(posedge clk)
    n231 <= infy_d1;
  /* fppowbf16.vhdl:5126:10  */
  always @(posedge clk)
    n232 <= s_nan_in;
  /* fppowbf16.vhdl:5126:10  */
  always @(posedge clk)
    n233 <= absxgtoneandnormal;
  /* fppowbf16.vhdl:5126:10  */
  always @(posedge clk)
    n234 <= absxgtoneandnormal_d1;
  /* fppowbf16.vhdl:5126:10  */
  always @(posedge clk)
    n235 <= absxltoneandnormal;
  /* fppowbf16.vhdl:5126:10  */
  always @(posedge clk)
    n236 <= absxltoneandnormal_d1;
  /* fppowbf16.vhdl:5126:10  */
  always @(posedge clk)
    n237 <= z_righty;
  /* fppowbf16.vhdl:5126:10  */
  always @(posedge clk)
    n238 <= weightlsbypre;
  /* fppowbf16.vhdl:5126:10  */
  always @(posedge clk)
    n239 <= weightlsby;
  /* fppowbf16.vhdl:5126:10  */
  always @(posedge clk)
    n240 <= oddinty;
endmodule

