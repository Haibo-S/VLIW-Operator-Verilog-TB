--------------------------------------------------------------------------------
--                  FixRealKCM_Freq500_uid8_T0_Freq500_uid11
-- VHDL generated for DummyFPGA @ 500MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 2
-- Target frequency (MHz): 500
-- Input signals: X
-- Output signals: Y
--  approx. input signal timings: X: (c0, 0.000000ns)
--  approx. output signal timings: Y: (c0, 0.550000ns)

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity FixRealKCM_Freq500_uid8_T0_Freq500_uid11 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(11 downto 0)   );
end entity;

architecture arch of FixRealKCM_Freq500_uid8_T0_Freq500_uid11 is
signal Y0 :  std_logic_vector(11 downto 0);
   -- timing of Y0: (c0, 0.550000ns)
signal Y1 :  std_logic_vector(11 downto 0);
   -- timing of Y1: (c0, 0.550000ns)
begin
   with X  select  Y0 <= 
      "000000001000" when "00000",
      "000001100100" when "00001",
      "000011000001" when "00010",
      "000100011101" when "00011",
      "000101111001" when "00100",
      "000111010110" when "00101",
      "001000110010" when "00110",
      "001010001110" when "00111",
      "001011101011" when "01000",
      "001101000111" when "01001",
      "001110100011" when "01010",
      "010000000000" when "01011",
      "010001011100" when "01100",
      "010010111000" when "01101",
      "010100010101" when "01110",
      "010101110001" when "01111",
      "010111001101" when "10000",
      "011000101010" when "10001",
      "011010000110" when "10010",
      "011011100010" when "10011",
      "011100111111" when "10100",
      "011110011011" when "10101",
      "011111110111" when "10110",
      "100001010100" when "10111",
      "100010110000" when "11000",
      "100100001100" when "11001",
      "100101101001" when "11010",
      "100111000101" when "11011",
      "101000100001" when "11100",
      "101001111110" when "11101",
      "101011011010" when "11110",
      "101100110110" when "11111",
      "------------" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                  FixRealKCM_Freq500_uid8_T1_Freq500_uid14
-- VHDL generated for DummyFPGA @ 500MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 2
-- Target frequency (MHz): 500
-- Input signals: X
-- Output signals: Y
--  approx. input signal timings: X: (c0, 0.000000ns)
--  approx. output signal timings: Y: (c0, 0.550000ns)

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity FixRealKCM_Freq500_uid8_T1_Freq500_uid14 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(6 downto 0)   );
end entity;

architecture arch of FixRealKCM_Freq500_uid8_T1_Freq500_uid14 is
signal Y0 :  std_logic_vector(6 downto 0);
   -- timing of Y0: (c0, 0.550000ns)
signal Y1 :  std_logic_vector(6 downto 0);
   -- timing of Y1: (c0, 0.550000ns)
begin
   with X  select  Y0 <= 
      "0000000" when "00000",
      "0000011" when "00001",
      "0000110" when "00010",
      "0001001" when "00011",
      "0001100" when "00100",
      "0001110" when "00101",
      "0010001" when "00110",
      "0010100" when "00111",
      "0010111" when "01000",
      "0011010" when "01001",
      "0011101" when "01010",
      "0100000" when "01011",
      "0100011" when "01100",
      "0100110" when "01101",
      "0101000" when "01110",
      "0101011" when "01111",
      "0101110" when "10000",
      "0110001" when "10001",
      "0110100" when "10010",
      "0110111" when "10011",
      "0111010" when "10100",
      "0111101" when "10101",
      "0111111" when "10110",
      "1000010" when "10111",
      "1000101" when "11000",
      "1001000" when "11001",
      "1001011" when "11010",
      "1001110" when "11011",
      "1010001" when "11100",
      "1010100" when "11101",
      "1010111" when "11110",
      "1011001" when "11111",
      "-------" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                 FixRealKCM_Freq500_uid20_T0_Freq500_uid23
-- VHDL generated for DummyFPGA @ 500MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 2
-- Target frequency (MHz): 500
-- Input signals: X
-- Output signals: Y
--  approx. input signal timings: X: (c0, 0.000000ns)
--  approx. output signal timings: Y: (c0, 0.550000ns)

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity FixRealKCM_Freq500_uid20_T0_Freq500_uid23 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(21 downto 0)   );
end entity;

architecture arch of FixRealKCM_Freq500_uid20_T0_Freq500_uid23 is
signal Y0 :  std_logic_vector(21 downto 0);
   -- timing of Y0: (c0, 0.550000ns)
signal Y1 :  std_logic_vector(21 downto 0);
   -- timing of Y1: (c0, 0.550000ns)
begin
   with X  select  Y0 <= 
      "0000000000000000000000" when "00000",
      "0000010110001011100100" when "00001",
      "0000101100010111001000" when "00010",
      "0001000010100010101101" when "00011",
      "0001011000101110010001" when "00100",
      "0001101110111001110101" when "00101",
      "0010000101000101011001" when "00110",
      "0010011011010000111101" when "00111",
      "0010110001011100100001" when "01000",
      "0011000111101000000110" when "01001",
      "0011011101110011101010" when "01010",
      "0011110011111111001110" when "01011",
      "0100001010001010110010" when "01100",
      "0100100000010110010110" when "01101",
      "0100110110100001111011" when "01110",
      "0101001100101101011111" when "01111",
      "0101100010111001000011" when "10000",
      "0101111001000100100111" when "10001",
      "0110001111010000001011" when "10010",
      "0110100101011011110000" when "10011",
      "0110111011100111010100" when "10100",
      "0111010001110010111000" when "10101",
      "0111100111111110011100" when "10110",
      "0111111110001010000000" when "10111",
      "1000010100010101100100" when "11000",
      "1000101010100001001001" when "11001",
      "1001000000101100101101" when "11010",
      "1001010110111000010001" when "11011",
      "1001101101000011110101" when "11100",
      "1010000011001111011001" when "11101",
      "1010011001011010111110" when "11110",
      "1010101111100110100010" when "11111",
      "----------------------" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                 FixRealKCM_Freq500_uid20_T1_Freq500_uid26
-- VHDL generated for DummyFPGA @ 500MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 2
-- Target frequency (MHz): 500
-- Input signals: X
-- Output signals: Y
--  approx. input signal timings: X: (c0, 0.000000ns)
--  approx. output signal timings: Y: (c0, 0.550000ns)

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity FixRealKCM_Freq500_uid20_T1_Freq500_uid26 is
    port (X : in  std_logic_vector(2 downto 0);
          Y : out  std_logic_vector(16 downto 0)   );
end entity;

architecture arch of FixRealKCM_Freq500_uid20_T1_Freq500_uid26 is
signal Y0 :  std_logic_vector(16 downto 0);
   -- timing of Y0: (c0, 0.550000ns)
signal Y1 :  std_logic_vector(16 downto 0);
   -- timing of Y1: (c0, 0.550000ns)
begin
   with X  select  Y0 <= 
      "00000000000000000" when "000",
      "00010110001011101" when "001",
      "00101100010111001" when "010",
      "01000010100010110" when "011",
      "01011000101110010" when "100",
      "01101110111001111" when "101",
      "10000101000101011" when "110",
      "10011011010001000" when "111",
      "-----------------" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                      FixFunctionByTable_Freq500_uid35
-- Evaluator for exp(x*1b-1) on [-1,1) for lsbIn=-9 (wIn=10), msbout=0, lsbOut=-14 (wOut=15). Out interval: [0.606531; 1.64711]. Output is unsigned

-- VHDL generated for DummyFPGA @ 500MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin (2010-2018)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 2
-- Target frequency (MHz): 500
-- Input signals: X
-- Output signals: Y
--  approx. input signal timings: X: (c0, 0.000000ns)
--  approx. output signal timings: Y: (c0, 0.550000ns)

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity FixFunctionByTable_Freq500_uid35 is
    port (X : in  std_logic_vector(9 downto 0);
          Y : out  std_logic_vector(14 downto 0)   );
end entity;

architecture arch of FixFunctionByTable_Freq500_uid35 is
signal Y0 :  std_logic_vector(14 downto 0);
   -- timing of Y0: (c0, 0.550000ns)
signal Y1 :  std_logic_vector(14 downto 0);
   -- timing of Y1: (c0, 0.550000ns)
begin
   with X  select  Y0 <= 
      "100000000000000" when "0000000000",
      "100000000010000" when "0000000001",
      "100000000100000" when "0000000010",
      "100000000110000" when "0000000011",
      "100000001000000" when "0000000100",
      "100000001010000" when "0000000101",
      "100000001100000" when "0000000110",
      "100000001110000" when "0000000111",
      "100000010000001" when "0000001000",
      "100000010010001" when "0000001001",
      "100000010100001" when "0000001010",
      "100000010110001" when "0000001011",
      "100000011000001" when "0000001100",
      "100000011010001" when "0000001101",
      "100000011100010" when "0000001110",
      "100000011110010" when "0000001111",
      "100000100000010" when "0000010000",
      "100000100010010" when "0000010001",
      "100000100100011" when "0000010010",
      "100000100110011" when "0000010011",
      "100000101000011" when "0000010100",
      "100000101010011" when "0000010101",
      "100000101100100" when "0000010110",
      "100000101110100" when "0000010111",
      "100000110000101" when "0000011000",
      "100000110010101" when "0000011001",
      "100000110100101" when "0000011010",
      "100000110110110" when "0000011011",
      "100000111000110" when "0000011100",
      "100000111010111" when "0000011101",
      "100000111100111" when "0000011110",
      "100000111111000" when "0000011111",
      "100001000001000" when "0000100000",
      "100001000011001" when "0000100001",
      "100001000101001" when "0000100010",
      "100001000111010" when "0000100011",
      "100001001001010" when "0000100100",
      "100001001011011" when "0000100101",
      "100001001101011" when "0000100110",
      "100001001111100" when "0000100111",
      "100001010001101" when "0000101000",
      "100001010011101" when "0000101001",
      "100001010101110" when "0000101010",
      "100001010111111" when "0000101011",
      "100001011001111" when "0000101100",
      "100001011100000" when "0000101101",
      "100001011110001" when "0000101110",
      "100001100000010" when "0000101111",
      "100001100010010" when "0000110000",
      "100001100100011" when "0000110001",
      "100001100110100" when "0000110010",
      "100001101000101" when "0000110011",
      "100001101010101" when "0000110100",
      "100001101100110" when "0000110101",
      "100001101110111" when "0000110110",
      "100001110001000" when "0000110111",
      "100001110011001" when "0000111000",
      "100001110101010" when "0000111001",
      "100001110111011" when "0000111010",
      "100001111001100" when "0000111011",
      "100001111011101" when "0000111100",
      "100001111101110" when "0000111101",
      "100001111111111" when "0000111110",
      "100010000010000" when "0000111111",
      "100010000100001" when "0001000000",
      "100010000110010" when "0001000001",
      "100010001000011" when "0001000010",
      "100010001010100" when "0001000011",
      "100010001100101" when "0001000100",
      "100010001110110" when "0001000101",
      "100010010000111" when "0001000110",
      "100010010011000" when "0001000111",
      "100010010101001" when "0001001000",
      "100010010111011" when "0001001001",
      "100010011001100" when "0001001010",
      "100010011011101" when "0001001011",
      "100010011101110" when "0001001100",
      "100010100000000" when "0001001101",
      "100010100010001" when "0001001110",
      "100010100100010" when "0001001111",
      "100010100110011" when "0001010000",
      "100010101000101" when "0001010001",
      "100010101010110" when "0001010010",
      "100010101100111" when "0001010011",
      "100010101111001" when "0001010100",
      "100010110001010" when "0001010101",
      "100010110011011" when "0001010110",
      "100010110101101" when "0001010111",
      "100010110111110" when "0001011000",
      "100010111010000" when "0001011001",
      "100010111100001" when "0001011010",
      "100010111110011" when "0001011011",
      "100011000000100" when "0001011100",
      "100011000010110" when "0001011101",
      "100011000100111" when "0001011110",
      "100011000111001" when "0001011111",
      "100011001001010" when "0001100000",
      "100011001011100" when "0001100001",
      "100011001101101" when "0001100010",
      "100011001111111" when "0001100011",
      "100011010010001" when "0001100100",
      "100011010100010" when "0001100101",
      "100011010110100" when "0001100110",
      "100011011000110" when "0001100111",
      "100011011010111" when "0001101000",
      "100011011101001" when "0001101001",
      "100011011111011" when "0001101010",
      "100011100001101" when "0001101011",
      "100011100011110" when "0001101100",
      "100011100110000" when "0001101101",
      "100011101000010" when "0001101110",
      "100011101010100" when "0001101111",
      "100011101100110" when "0001110000",
      "100011101111000" when "0001110001",
      "100011110001001" when "0001110010",
      "100011110011011" when "0001110011",
      "100011110101101" when "0001110100",
      "100011110111111" when "0001110101",
      "100011111010001" when "0001110110",
      "100011111100011" when "0001110111",
      "100011111110101" when "0001111000",
      "100100000000111" when "0001111001",
      "100100000011001" when "0001111010",
      "100100000101011" when "0001111011",
      "100100000111101" when "0001111100",
      "100100001001111" when "0001111101",
      "100100001100001" when "0001111110",
      "100100001110011" when "0001111111",
      "100100010000110" when "0010000000",
      "100100010011000" when "0010000001",
      "100100010101010" when "0010000010",
      "100100010111100" when "0010000011",
      "100100011001110" when "0010000100",
      "100100011100000" when "0010000101",
      "100100011110011" when "0010000110",
      "100100100000101" when "0010000111",
      "100100100010111" when "0010001000",
      "100100100101001" when "0010001001",
      "100100100111100" when "0010001010",
      "100100101001110" when "0010001011",
      "100100101100000" when "0010001100",
      "100100101110011" when "0010001101",
      "100100110000101" when "0010001110",
      "100100110010111" when "0010001111",
      "100100110101010" when "0010010000",
      "100100110111100" when "0010010001",
      "100100111001111" when "0010010010",
      "100100111100001" when "0010010011",
      "100100111110100" when "0010010100",
      "100101000000110" when "0010010101",
      "100101000011001" when "0010010110",
      "100101000101011" when "0010010111",
      "100101000111110" when "0010011000",
      "100101001010000" when "0010011001",
      "100101001100011" when "0010011010",
      "100101001110110" when "0010011011",
      "100101010001000" when "0010011100",
      "100101010011011" when "0010011101",
      "100101010101101" when "0010011110",
      "100101011000000" when "0010011111",
      "100101011010011" when "0010100000",
      "100101011100110" when "0010100001",
      "100101011111000" when "0010100010",
      "100101100001011" when "0010100011",
      "100101100011110" when "0010100100",
      "100101100110001" when "0010100101",
      "100101101000011" when "0010100110",
      "100101101010110" when "0010100111",
      "100101101101001" when "0010101000",
      "100101101111100" when "0010101001",
      "100101110001111" when "0010101010",
      "100101110100010" when "0010101011",
      "100101110110101" when "0010101100",
      "100101111001000" when "0010101101",
      "100101111011011" when "0010101110",
      "100101111101101" when "0010101111",
      "100110000000000" when "0010110000",
      "100110000010011" when "0010110001",
      "100110000100111" when "0010110010",
      "100110000111010" when "0010110011",
      "100110001001101" when "0010110100",
      "100110001100000" when "0010110101",
      "100110001110011" when "0010110110",
      "100110010000110" when "0010110111",
      "100110010011001" when "0010111000",
      "100110010101100" when "0010111001",
      "100110010111111" when "0010111010",
      "100110011010011" when "0010111011",
      "100110011100110" when "0010111100",
      "100110011111001" when "0010111101",
      "100110100001100" when "0010111110",
      "100110100100000" when "0010111111",
      "100110100110011" when "0011000000",
      "100110101000110" when "0011000001",
      "100110101011010" when "0011000010",
      "100110101101101" when "0011000011",
      "100110110000000" when "0011000100",
      "100110110010100" when "0011000101",
      "100110110100111" when "0011000110",
      "100110110111010" when "0011000111",
      "100110111001110" when "0011001000",
      "100110111100001" when "0011001001",
      "100110111110101" when "0011001010",
      "100111000001000" when "0011001011",
      "100111000011100" when "0011001100",
      "100111000101111" when "0011001101",
      "100111001000011" when "0011001110",
      "100111001010111" when "0011001111",
      "100111001101010" when "0011010000",
      "100111001111110" when "0011010001",
      "100111010010001" when "0011010010",
      "100111010100101" when "0011010011",
      "100111010111001" when "0011010100",
      "100111011001100" when "0011010101",
      "100111011100000" when "0011010110",
      "100111011110100" when "0011010111",
      "100111100001000" when "0011011000",
      "100111100011011" when "0011011001",
      "100111100101111" when "0011011010",
      "100111101000011" when "0011011011",
      "100111101010111" when "0011011100",
      "100111101101011" when "0011011101",
      "100111101111110" when "0011011110",
      "100111110010010" when "0011011111",
      "100111110100110" when "0011100000",
      "100111110111010" when "0011100001",
      "100111111001110" when "0011100010",
      "100111111100010" when "0011100011",
      "100111111110110" when "0011100100",
      "101000000001010" when "0011100101",
      "101000000011110" when "0011100110",
      "101000000110010" when "0011100111",
      "101000001000110" when "0011101000",
      "101000001011010" when "0011101001",
      "101000001101110" when "0011101010",
      "101000010000010" when "0011101011",
      "101000010010111" when "0011101100",
      "101000010101011" when "0011101101",
      "101000010111111" when "0011101110",
      "101000011010011" when "0011101111",
      "101000011100111" when "0011110000",
      "101000011111100" when "0011110001",
      "101000100010000" when "0011110010",
      "101000100100100" when "0011110011",
      "101000100111000" when "0011110100",
      "101000101001101" when "0011110101",
      "101000101100001" when "0011110110",
      "101000101110101" when "0011110111",
      "101000110001010" when "0011111000",
      "101000110011110" when "0011111001",
      "101000110110011" when "0011111010",
      "101000111000111" when "0011111011",
      "101000111011011" when "0011111100",
      "101000111110000" when "0011111101",
      "101001000000100" when "0011111110",
      "101001000011001" when "0011111111",
      "101001000101101" when "0100000000",
      "101001001000010" when "0100000001",
      "101001001010111" when "0100000010",
      "101001001101011" when "0100000011",
      "101001010000000" when "0100000100",
      "101001010010100" when "0100000101",
      "101001010101001" when "0100000110",
      "101001010111110" when "0100000111",
      "101001011010010" when "0100001000",
      "101001011100111" when "0100001001",
      "101001011111100" when "0100001010",
      "101001100010001" when "0100001011",
      "101001100100101" when "0100001100",
      "101001100111010" when "0100001101",
      "101001101001111" when "0100001110",
      "101001101100100" when "0100001111",
      "101001101111001" when "0100010000",
      "101001110001110" when "0100010001",
      "101001110100011" when "0100010010",
      "101001110110111" when "0100010011",
      "101001111001100" when "0100010100",
      "101001111100001" when "0100010101",
      "101001111110110" when "0100010110",
      "101010000001011" when "0100010111",
      "101010000100000" when "0100011000",
      "101010000110101" when "0100011001",
      "101010001001010" when "0100011010",
      "101010001100000" when "0100011011",
      "101010001110101" when "0100011100",
      "101010010001010" when "0100011101",
      "101010010011111" when "0100011110",
      "101010010110100" when "0100011111",
      "101010011001001" when "0100100000",
      "101010011011110" when "0100100001",
      "101010011110100" when "0100100010",
      "101010100001001" when "0100100011",
      "101010100011110" when "0100100100",
      "101010100110100" when "0100100101",
      "101010101001001" when "0100100110",
      "101010101011110" when "0100100111",
      "101010101110100" when "0100101000",
      "101010110001001" when "0100101001",
      "101010110011110" when "0100101010",
      "101010110110100" when "0100101011",
      "101010111001001" when "0100101100",
      "101010111011111" when "0100101101",
      "101010111110100" when "0100101110",
      "101011000001010" when "0100101111",
      "101011000011111" when "0100110000",
      "101011000110101" when "0100110001",
      "101011001001010" when "0100110010",
      "101011001100000" when "0100110011",
      "101011001110101" when "0100110100",
      "101011010001011" when "0100110101",
      "101011010100001" when "0100110110",
      "101011010110110" when "0100110111",
      "101011011001100" when "0100111000",
      "101011011100010" when "0100111001",
      "101011011110111" when "0100111010",
      "101011100001101" when "0100111011",
      "101011100100011" when "0100111100",
      "101011100111001" when "0100111101",
      "101011101001111" when "0100111110",
      "101011101100100" when "0100111111",
      "101011101111010" when "0101000000",
      "101011110010000" when "0101000001",
      "101011110100110" when "0101000010",
      "101011110111100" when "0101000011",
      "101011111010010" when "0101000100",
      "101011111101000" when "0101000101",
      "101011111111110" when "0101000110",
      "101100000010100" when "0101000111",
      "101100000101010" when "0101001000",
      "101100001000000" when "0101001001",
      "101100001010110" when "0101001010",
      "101100001101100" when "0101001011",
      "101100010000010" when "0101001100",
      "101100010011000" when "0101001101",
      "101100010101111" when "0101001110",
      "101100011000101" when "0101001111",
      "101100011011011" when "0101010000",
      "101100011110001" when "0101010001",
      "101100100000111" when "0101010010",
      "101100100011110" when "0101010011",
      "101100100110100" when "0101010100",
      "101100101001010" when "0101010101",
      "101100101100001" when "0101010110",
      "101100101110111" when "0101010111",
      "101100110001101" when "0101011000",
      "101100110100100" when "0101011001",
      "101100110111010" when "0101011010",
      "101100111010001" when "0101011011",
      "101100111100111" when "0101011100",
      "101100111111110" when "0101011101",
      "101101000010100" when "0101011110",
      "101101000101011" when "0101011111",
      "101101001000001" when "0101100000",
      "101101001011000" when "0101100001",
      "101101001101110" when "0101100010",
      "101101010000101" when "0101100011",
      "101101010011100" when "0101100100",
      "101101010110010" when "0101100101",
      "101101011001001" when "0101100110",
      "101101011100000" when "0101100111",
      "101101011110110" when "0101101000",
      "101101100001101" when "0101101001",
      "101101100100100" when "0101101010",
      "101101100111011" when "0101101011",
      "101101101010001" when "0101101100",
      "101101101101000" when "0101101101",
      "101101101111111" when "0101101110",
      "101101110010110" when "0101101111",
      "101101110101101" when "0101110000",
      "101101111000100" when "0101110001",
      "101101111011011" when "0101110010",
      "101101111110010" when "0101110011",
      "101110000001001" when "0101110100",
      "101110000100000" when "0101110101",
      "101110000110111" when "0101110110",
      "101110001001110" when "0101110111",
      "101110001100101" when "0101111000",
      "101110001111100" when "0101111001",
      "101110010010011" when "0101111010",
      "101110010101010" when "0101111011",
      "101110011000010" when "0101111100",
      "101110011011001" when "0101111101",
      "101110011110000" when "0101111110",
      "101110100000111" when "0101111111",
      "101110100011111" when "0110000000",
      "101110100110110" when "0110000001",
      "101110101001101" when "0110000010",
      "101110101100101" when "0110000011",
      "101110101111100" when "0110000100",
      "101110110010011" when "0110000101",
      "101110110101011" when "0110000110",
      "101110111000010" when "0110000111",
      "101110111011010" when "0110001000",
      "101110111110001" when "0110001001",
      "101111000001001" when "0110001010",
      "101111000100000" when "0110001011",
      "101111000111000" when "0110001100",
      "101111001001111" when "0110001101",
      "101111001100111" when "0110001110",
      "101111001111110" when "0110001111",
      "101111010010110" when "0110010000",
      "101111010101110" when "0110010001",
      "101111011000101" when "0110010010",
      "101111011011101" when "0110010011",
      "101111011110101" when "0110010100",
      "101111100001101" when "0110010101",
      "101111100100100" when "0110010110",
      "101111100111100" when "0110010111",
      "101111101010100" when "0110011000",
      "101111101101100" when "0110011001",
      "101111110000100" when "0110011010",
      "101111110011011" when "0110011011",
      "101111110110011" when "0110011100",
      "101111111001011" when "0110011101",
      "101111111100011" when "0110011110",
      "101111111111011" when "0110011111",
      "110000000010011" when "0110100000",
      "110000000101011" when "0110100001",
      "110000001000011" when "0110100010",
      "110000001011011" when "0110100011",
      "110000001110100" when "0110100100",
      "110000010001100" when "0110100101",
      "110000010100100" when "0110100110",
      "110000010111100" when "0110100111",
      "110000011010100" when "0110101000",
      "110000011101100" when "0110101001",
      "110000100000101" when "0110101010",
      "110000100011101" when "0110101011",
      "110000100110101" when "0110101100",
      "110000101001110" when "0110101101",
      "110000101100110" when "0110101110",
      "110000101111110" when "0110101111",
      "110000110010111" when "0110110000",
      "110000110101111" when "0110110001",
      "110000111000111" when "0110110010",
      "110000111100000" when "0110110011",
      "110000111111000" when "0110110100",
      "110001000010001" when "0110110101",
      "110001000101001" when "0110110110",
      "110001001000010" when "0110110111",
      "110001001011011" when "0110111000",
      "110001001110011" when "0110111001",
      "110001010001100" when "0110111010",
      "110001010100100" when "0110111011",
      "110001010111101" when "0110111100",
      "110001011010110" when "0110111101",
      "110001011101111" when "0110111110",
      "110001100000111" when "0110111111",
      "110001100100000" when "0111000000",
      "110001100111001" when "0111000001",
      "110001101010010" when "0111000010",
      "110001101101010" when "0111000011",
      "110001110000011" when "0111000100",
      "110001110011100" when "0111000101",
      "110001110110101" when "0111000110",
      "110001111001110" when "0111000111",
      "110001111100111" when "0111001000",
      "110010000000000" when "0111001001",
      "110010000011001" when "0111001010",
      "110010000110010" when "0111001011",
      "110010001001011" when "0111001100",
      "110010001100100" when "0111001101",
      "110010001111101" when "0111001110",
      "110010010010110" when "0111001111",
      "110010010110000" when "0111010000",
      "110010011001001" when "0111010001",
      "110010011100010" when "0111010010",
      "110010011111011" when "0111010011",
      "110010100010101" when "0111010100",
      "110010100101110" when "0111010101",
      "110010101000111" when "0111010110",
      "110010101100000" when "0111010111",
      "110010101111010" when "0111011000",
      "110010110010011" when "0111011001",
      "110010110101101" when "0111011010",
      "110010111000110" when "0111011011",
      "110010111011111" when "0111011100",
      "110010111111001" when "0111011101",
      "110011000010010" when "0111011110",
      "110011000101100" when "0111011111",
      "110011001000110" when "0111100000",
      "110011001011111" when "0111100001",
      "110011001111001" when "0111100010",
      "110011010010010" when "0111100011",
      "110011010101100" when "0111100100",
      "110011011000110" when "0111100101",
      "110011011011111" when "0111100110",
      "110011011111001" when "0111100111",
      "110011100010011" when "0111101000",
      "110011100101101" when "0111101001",
      "110011101000110" when "0111101010",
      "110011101100000" when "0111101011",
      "110011101111010" when "0111101100",
      "110011110010100" when "0111101101",
      "110011110101110" when "0111101110",
      "110011111001000" when "0111101111",
      "110011111100010" when "0111110000",
      "110011111111100" when "0111110001",
      "110100000010110" when "0111110010",
      "110100000110000" when "0111110011",
      "110100001001010" when "0111110100",
      "110100001100100" when "0111110101",
      "110100001111110" when "0111110110",
      "110100010011000" when "0111110111",
      "110100010110010" when "0111111000",
      "110100011001101" when "0111111001",
      "110100011100111" when "0111111010",
      "110100100000001" when "0111111011",
      "110100100011011" when "0111111100",
      "110100100110110" when "0111111101",
      "110100101010000" when "0111111110",
      "110100101101010" when "0111111111",
      "010011011010001" when "1000000000",
      "010011011011011" when "1000000001",
      "010011011100101" when "1000000010",
      "010011011101111" when "1000000011",
      "010011011111000" when "1000000100",
      "010011100000010" when "1000000101",
      "010011100001100" when "1000000110",
      "010011100010110" when "1000000111",
      "010011100011111" when "1000001000",
      "010011100101001" when "1000001001",
      "010011100110011" when "1000001010",
      "010011100111101" when "1000001011",
      "010011101000111" when "1000001100",
      "010011101010000" when "1000001101",
      "010011101011010" when "1000001110",
      "010011101100100" when "1000001111",
      "010011101101110" when "1000010000",
      "010011101111000" when "1000010001",
      "010011110000010" when "1000010010",
      "010011110001100" when "1000010011",
      "010011110010101" when "1000010100",
      "010011110011111" when "1000010101",
      "010011110101001" when "1000010110",
      "010011110110011" when "1000010111",
      "010011110111101" when "1000011000",
      "010011111000111" when "1000011001",
      "010011111010001" when "1000011010",
      "010011111011011" when "1000011011",
      "010011111100101" when "1000011100",
      "010011111101111" when "1000011101",
      "010011111111001" when "1000011110",
      "010100000000011" when "1000011111",
      "010100000001101" when "1000100000",
      "010100000010111" when "1000100001",
      "010100000100001" when "1000100010",
      "010100000101011" when "1000100011",
      "010100000110101" when "1000100100",
      "010100000111111" when "1000100101",
      "010100001001001" when "1000100110",
      "010100001010011" when "1000100111",
      "010100001011101" when "1000101000",
      "010100001100111" when "1000101001",
      "010100001110001" when "1000101010",
      "010100001111100" when "1000101011",
      "010100010000110" when "1000101100",
      "010100010010000" when "1000101101",
      "010100010011010" when "1000101110",
      "010100010100100" when "1000101111",
      "010100010101110" when "1000110000",
      "010100010111000" when "1000110001",
      "010100011000011" when "1000110010",
      "010100011001101" when "1000110011",
      "010100011010111" when "1000110100",
      "010100011100001" when "1000110101",
      "010100011101100" when "1000110110",
      "010100011110110" when "1000110111",
      "010100100000000" when "1000111000",
      "010100100001010" when "1000111001",
      "010100100010101" when "1000111010",
      "010100100011111" when "1000111011",
      "010100100101001" when "1000111100",
      "010100100110011" when "1000111101",
      "010100100111110" when "1000111110",
      "010100101001000" when "1000111111",
      "010100101010010" when "1001000000",
      "010100101011101" when "1001000001",
      "010100101100111" when "1001000010",
      "010100101110001" when "1001000011",
      "010100101111100" when "1001000100",
      "010100110000110" when "1001000101",
      "010100110010000" when "1001000110",
      "010100110011011" when "1001000111",
      "010100110100101" when "1001001000",
      "010100110110000" when "1001001001",
      "010100110111010" when "1001001010",
      "010100111000101" when "1001001011",
      "010100111001111" when "1001001100",
      "010100111011001" when "1001001101",
      "010100111100100" when "1001001110",
      "010100111101110" when "1001001111",
      "010100111111001" when "1001010000",
      "010101000000011" when "1001010001",
      "010101000001110" when "1001010010",
      "010101000011000" when "1001010011",
      "010101000100011" when "1001010100",
      "010101000101101" when "1001010101",
      "010101000111000" when "1001010110",
      "010101001000011" when "1001010111",
      "010101001001101" when "1001011000",
      "010101001011000" when "1001011001",
      "010101001100010" when "1001011010",
      "010101001101101" when "1001011011",
      "010101001111000" when "1001011100",
      "010101010000010" when "1001011101",
      "010101010001101" when "1001011110",
      "010101010010111" when "1001011111",
      "010101010100010" when "1001100000",
      "010101010101101" when "1001100001",
      "010101010110111" when "1001100010",
      "010101011000010" when "1001100011",
      "010101011001101" when "1001100100",
      "010101011011000" when "1001100101",
      "010101011100010" when "1001100110",
      "010101011101101" when "1001100111",
      "010101011111000" when "1001101000",
      "010101100000010" when "1001101001",
      "010101100001101" when "1001101010",
      "010101100011000" when "1001101011",
      "010101100100011" when "1001101100",
      "010101100101110" when "1001101101",
      "010101100111000" when "1001101110",
      "010101101000011" when "1001101111",
      "010101101001110" when "1001110000",
      "010101101011001" when "1001110001",
      "010101101100100" when "1001110010",
      "010101101101110" when "1001110011",
      "010101101111001" when "1001110100",
      "010101110000100" when "1001110101",
      "010101110001111" when "1001110110",
      "010101110011010" when "1001110111",
      "010101110100101" when "1001111000",
      "010101110110000" when "1001111001",
      "010101110111011" when "1001111010",
      "010101111000110" when "1001111011",
      "010101111010001" when "1001111100",
      "010101111011100" when "1001111101",
      "010101111100111" when "1001111110",
      "010101111110010" when "1001111111",
      "010101111111101" when "1010000000",
      "010110000001000" when "1010000001",
      "010110000010011" when "1010000010",
      "010110000011110" when "1010000011",
      "010110000101001" when "1010000100",
      "010110000110100" when "1010000101",
      "010110000111111" when "1010000110",
      "010110001001010" when "1010000111",
      "010110001010101" when "1010001000",
      "010110001100000" when "1010001001",
      "010110001101011" when "1010001010",
      "010110001110110" when "1010001011",
      "010110010000001" when "1010001100",
      "010110010001100" when "1010001101",
      "010110010011000" when "1010001110",
      "010110010100011" when "1010001111",
      "010110010101110" when "1010010000",
      "010110010111001" when "1010010001",
      "010110011000100" when "1010010010",
      "010110011001111" when "1010010011",
      "010110011011011" when "1010010100",
      "010110011100110" when "1010010101",
      "010110011110001" when "1010010110",
      "010110011111100" when "1010010111",
      "010110100001000" when "1010011000",
      "010110100010011" when "1010011001",
      "010110100011110" when "1010011010",
      "010110100101001" when "1010011011",
      "010110100110101" when "1010011100",
      "010110101000000" when "1010011101",
      "010110101001011" when "1010011110",
      "010110101010111" when "1010011111",
      "010110101100010" when "1010100000",
      "010110101101101" when "1010100001",
      "010110101111001" when "1010100010",
      "010110110000100" when "1010100011",
      "010110110001111" when "1010100100",
      "010110110011011" when "1010100101",
      "010110110100110" when "1010100110",
      "010110110110010" when "1010100111",
      "010110110111101" when "1010101000",
      "010110111001001" when "1010101001",
      "010110111010100" when "1010101010",
      "010110111011111" when "1010101011",
      "010110111101011" when "1010101100",
      "010110111110110" when "1010101101",
      "010111000000010" when "1010101110",
      "010111000001101" when "1010101111",
      "010111000011001" when "1010110000",
      "010111000100100" when "1010110001",
      "010111000110000" when "1010110010",
      "010111000111100" when "1010110011",
      "010111001000111" when "1010110100",
      "010111001010011" when "1010110101",
      "010111001011110" when "1010110110",
      "010111001101010" when "1010110111",
      "010111001110110" when "1010111000",
      "010111010000001" when "1010111001",
      "010111010001101" when "1010111010",
      "010111010011000" when "1010111011",
      "010111010100100" when "1010111100",
      "010111010110000" when "1010111101",
      "010111010111011" when "1010111110",
      "010111011000111" when "1010111111",
      "010111011010011" when "1011000000",
      "010111011011111" when "1011000001",
      "010111011101010" when "1011000010",
      "010111011110110" when "1011000011",
      "010111100000010" when "1011000100",
      "010111100001101" when "1011000101",
      "010111100011001" when "1011000110",
      "010111100100101" when "1011000111",
      "010111100110001" when "1011001000",
      "010111100111101" when "1011001001",
      "010111101001000" when "1011001010",
      "010111101010100" when "1011001011",
      "010111101100000" when "1011001100",
      "010111101101100" when "1011001101",
      "010111101111000" when "1011001110",
      "010111110000100" when "1011001111",
      "010111110010000" when "1011010000",
      "010111110011011" when "1011010001",
      "010111110100111" when "1011010010",
      "010111110110011" when "1011010011",
      "010111110111111" when "1011010100",
      "010111111001011" when "1011010101",
      "010111111010111" when "1011010110",
      "010111111100011" when "1011010111",
      "010111111101111" when "1011011000",
      "010111111111011" when "1011011001",
      "011000000000111" when "1011011010",
      "011000000010011" when "1011011011",
      "011000000011111" when "1011011100",
      "011000000101011" when "1011011101",
      "011000000110111" when "1011011110",
      "011000001000011" when "1011011111",
      "011000001001111" when "1011100000",
      "011000001011011" when "1011100001",
      "011000001100111" when "1011100010",
      "011000001110100" when "1011100011",
      "011000010000000" when "1011100100",
      "011000010001100" when "1011100101",
      "011000010011000" when "1011100110",
      "011000010100100" when "1011100111",
      "011000010110000" when "1011101000",
      "011000010111100" when "1011101001",
      "011000011001001" when "1011101010",
      "011000011010101" when "1011101011",
      "011000011100001" when "1011101100",
      "011000011101101" when "1011101101",
      "011000011111010" when "1011101110",
      "011000100000110" when "1011101111",
      "011000100010010" when "1011110000",
      "011000100011110" when "1011110001",
      "011000100101011" when "1011110010",
      "011000100110111" when "1011110011",
      "011000101000011" when "1011110100",
      "011000101010000" when "1011110101",
      "011000101011100" when "1011110110",
      "011000101101000" when "1011110111",
      "011000101110101" when "1011111000",
      "011000110000001" when "1011111001",
      "011000110001101" when "1011111010",
      "011000110011010" when "1011111011",
      "011000110100110" when "1011111100",
      "011000110110011" when "1011111101",
      "011000110111111" when "1011111110",
      "011000111001011" when "1011111111",
      "011000111011000" when "1100000000",
      "011000111100100" when "1100000001",
      "011000111110001" when "1100000010",
      "011000111111101" when "1100000011",
      "011001000001010" when "1100000100",
      "011001000010110" when "1100000101",
      "011001000100011" when "1100000110",
      "011001000101111" when "1100000111",
      "011001000111100" when "1100001000",
      "011001001001001" when "1100001001",
      "011001001010101" when "1100001010",
      "011001001100010" when "1100001011",
      "011001001101110" when "1100001100",
      "011001001111011" when "1100001101",
      "011001010001000" when "1100001110",
      "011001010010100" when "1100001111",
      "011001010100001" when "1100010000",
      "011001010101101" when "1100010001",
      "011001010111010" when "1100010010",
      "011001011000111" when "1100010011",
      "011001011010100" when "1100010100",
      "011001011100000" when "1100010101",
      "011001011101101" when "1100010110",
      "011001011111010" when "1100010111",
      "011001100000110" when "1100011000",
      "011001100010011" when "1100011001",
      "011001100100000" when "1100011010",
      "011001100101101" when "1100011011",
      "011001100111010" when "1100011100",
      "011001101000110" when "1100011101",
      "011001101010011" when "1100011110",
      "011001101100000" when "1100011111",
      "011001101101101" when "1100100000",
      "011001101111010" when "1100100001",
      "011001110000111" when "1100100010",
      "011001110010100" when "1100100011",
      "011001110100000" when "1100100100",
      "011001110101101" when "1100100101",
      "011001110111010" when "1100100110",
      "011001111000111" when "1100100111",
      "011001111010100" when "1100101000",
      "011001111100001" when "1100101001",
      "011001111101110" when "1100101010",
      "011001111111011" when "1100101011",
      "011010000001000" when "1100101100",
      "011010000010101" when "1100101101",
      "011010000100010" when "1100101110",
      "011010000101111" when "1100101111",
      "011010000111100" when "1100110000",
      "011010001001001" when "1100110001",
      "011010001010110" when "1100110010",
      "011010001100011" when "1100110011",
      "011010001110001" when "1100110100",
      "011010001111110" when "1100110101",
      "011010010001011" when "1100110110",
      "011010010011000" when "1100110111",
      "011010010100101" when "1100111000",
      "011010010110010" when "1100111001",
      "011010010111111" when "1100111010",
      "011010011001101" when "1100111011",
      "011010011011010" when "1100111100",
      "011010011100111" when "1100111101",
      "011010011110100" when "1100111110",
      "011010100000010" when "1100111111",
      "011010100001111" when "1101000000",
      "011010100011100" when "1101000001",
      "011010100101001" when "1101000010",
      "011010100110111" when "1101000011",
      "011010101000100" when "1101000100",
      "011010101010001" when "1101000101",
      "011010101011111" when "1101000110",
      "011010101101100" when "1101000111",
      "011010101111001" when "1101001000",
      "011010110000111" when "1101001001",
      "011010110010100" when "1101001010",
      "011010110100010" when "1101001011",
      "011010110101111" when "1101001100",
      "011010110111100" when "1101001101",
      "011010111001010" when "1101001110",
      "011010111010111" when "1101001111",
      "011010111100101" when "1101010000",
      "011010111110010" when "1101010001",
      "011011000000000" when "1101010010",
      "011011000001101" when "1101010011",
      "011011000011011" when "1101010100",
      "011011000101000" when "1101010101",
      "011011000110110" when "1101010110",
      "011011001000011" when "1101010111",
      "011011001010001" when "1101011000",
      "011011001011111" when "1101011001",
      "011011001101100" when "1101011010",
      "011011001111010" when "1101011011",
      "011011010000111" when "1101011100",
      "011011010010101" when "1101011101",
      "011011010100011" when "1101011110",
      "011011010110000" when "1101011111",
      "011011010111110" when "1101100000",
      "011011011001100" when "1101100001",
      "011011011011001" when "1101100010",
      "011011011100111" when "1101100011",
      "011011011110101" when "1101100100",
      "011011100000011" when "1101100101",
      "011011100010000" when "1101100110",
      "011011100011110" when "1101100111",
      "011011100101100" when "1101101000",
      "011011100111010" when "1101101001",
      "011011101001000" when "1101101010",
      "011011101010101" when "1101101011",
      "011011101100011" when "1101101100",
      "011011101110001" when "1101101101",
      "011011101111111" when "1101101110",
      "011011110001101" when "1101101111",
      "011011110011011" when "1101110000",
      "011011110101001" when "1101110001",
      "011011110110110" when "1101110010",
      "011011111000100" when "1101110011",
      "011011111010010" when "1101110100",
      "011011111100000" when "1101110101",
      "011011111101110" when "1101110110",
      "011011111111100" when "1101110111",
      "011100000001010" when "1101111000",
      "011100000011000" when "1101111001",
      "011100000100110" when "1101111010",
      "011100000110100" when "1101111011",
      "011100001000010" when "1101111100",
      "011100001010001" when "1101111101",
      "011100001011111" when "1101111110",
      "011100001101101" when "1101111111",
      "011100001111011" when "1110000000",
      "011100010001001" when "1110000001",
      "011100010010111" when "1110000010",
      "011100010100101" when "1110000011",
      "011100010110011" when "1110000100",
      "011100011000010" when "1110000101",
      "011100011010000" when "1110000110",
      "011100011011110" when "1110000111",
      "011100011101100" when "1110001000",
      "011100011111010" when "1110001001",
      "011100100001001" when "1110001010",
      "011100100010111" when "1110001011",
      "011100100100101" when "1110001100",
      "011100100110100" when "1110001101",
      "011100101000010" when "1110001110",
      "011100101010000" when "1110001111",
      "011100101011111" when "1110010000",
      "011100101101101" when "1110010001",
      "011100101111011" when "1110010010",
      "011100110001010" when "1110010011",
      "011100110011000" when "1110010100",
      "011100110100110" when "1110010101",
      "011100110110101" when "1110010110",
      "011100111000011" when "1110010111",
      "011100111010010" when "1110011000",
      "011100111100000" when "1110011001",
      "011100111101111" when "1110011010",
      "011100111111101" when "1110011011",
      "011101000001100" when "1110011100",
      "011101000011010" when "1110011101",
      "011101000101001" when "1110011110",
      "011101000110111" when "1110011111",
      "011101001000110" when "1110100000",
      "011101001010100" when "1110100001",
      "011101001100011" when "1110100010",
      "011101001110010" when "1110100011",
      "011101010000000" when "1110100100",
      "011101010001111" when "1110100101",
      "011101010011101" when "1110100110",
      "011101010101100" when "1110100111",
      "011101010111011" when "1110101000",
      "011101011001001" when "1110101001",
      "011101011011000" when "1110101010",
      "011101011100111" when "1110101011",
      "011101011110110" when "1110101100",
      "011101100000100" when "1110101101",
      "011101100010011" when "1110101110",
      "011101100100010" when "1110101111",
      "011101100110001" when "1110110000",
      "011101101000000" when "1110110001",
      "011101101001110" when "1110110010",
      "011101101011101" when "1110110011",
      "011101101101100" when "1110110100",
      "011101101111011" when "1110110101",
      "011101110001010" when "1110110110",
      "011101110011001" when "1110110111",
      "011101110101000" when "1110111000",
      "011101110110110" when "1110111001",
      "011101111000101" when "1110111010",
      "011101111010100" when "1110111011",
      "011101111100011" when "1110111100",
      "011101111110010" when "1110111101",
      "011110000000001" when "1110111110",
      "011110000010000" when "1110111111",
      "011110000011111" when "1111000000",
      "011110000101110" when "1111000001",
      "011110000111101" when "1111000010",
      "011110001001101" when "1111000011",
      "011110001011100" when "1111000100",
      "011110001101011" when "1111000101",
      "011110001111010" when "1111000110",
      "011110010001001" when "1111000111",
      "011110010011000" when "1111001000",
      "011110010100111" when "1111001001",
      "011110010110110" when "1111001010",
      "011110011000110" when "1111001011",
      "011110011010101" when "1111001100",
      "011110011100100" when "1111001101",
      "011110011110011" when "1111001110",
      "011110100000010" when "1111001111",
      "011110100010010" when "1111010000",
      "011110100100001" when "1111010001",
      "011110100110000" when "1111010010",
      "011110101000000" when "1111010011",
      "011110101001111" when "1111010100",
      "011110101011110" when "1111010101",
      "011110101101110" when "1111010110",
      "011110101111101" when "1111010111",
      "011110110001100" when "1111011000",
      "011110110011100" when "1111011001",
      "011110110101011" when "1111011010",
      "011110110111011" when "1111011011",
      "011110111001010" when "1111011100",
      "011110111011001" when "1111011101",
      "011110111101001" when "1111011110",
      "011110111111000" when "1111011111",
      "011111000001000" when "1111100000",
      "011111000010111" when "1111100001",
      "011111000100111" when "1111100010",
      "011111000110111" when "1111100011",
      "011111001000110" when "1111100100",
      "011111001010110" when "1111100101",
      "011111001100101" when "1111100110",
      "011111001110101" when "1111100111",
      "011111010000100" when "1111101000",
      "011111010010100" when "1111101001",
      "011111010100100" when "1111101010",
      "011111010110011" when "1111101011",
      "011111011000011" when "1111101100",
      "011111011010011" when "1111101101",
      "011111011100011" when "1111101110",
      "011111011110010" when "1111101111",
      "011111100000010" when "1111110000",
      "011111100010010" when "1111110001",
      "011111100100010" when "1111110010",
      "011111100110001" when "1111110011",
      "011111101000001" when "1111110100",
      "011111101010001" when "1111110101",
      "011111101100001" when "1111110110",
      "011111101110001" when "1111110111",
      "011111110000000" when "1111111000",
      "011111110010000" when "1111111001",
      "011111110100000" when "1111111010",
      "011111110110000" when "1111111011",
      "011111111000000" when "1111111100",
      "011111111010000" when "1111111101",
      "011111111100000" when "1111111110",
      "011111111110000" when "1111111111",
      "---------------" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                      FixFunctionByTable_Freq500_uid38
-- Evaluator for (exp(x*1b-11)-1) on [-1,1) for lsbIn=-3 (wIn=4), msbout=-11, lsbOut=-14 (wOut=4). Out interval: [-0.000488162; 0.000427337]. Output is signed

-- VHDL generated for DummyFPGA @ 500MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin (2010-2018)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 2
-- Target frequency (MHz): 500
-- Input signals: X
-- Output signals: Y
--  approx. input signal timings: X: (c0, 0.000000ns)
--  approx. output signal timings: Y: (c0, 0.550000ns)

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity FixFunctionByTable_Freq500_uid38 is
    port (X : in  std_logic_vector(3 downto 0);
          Y : out  std_logic_vector(3 downto 0)   );
end entity;

architecture arch of FixFunctionByTable_Freq500_uid38 is
signal Y0 :  std_logic_vector(3 downto 0);
   -- timing of Y0: (c0, 0.550000ns)
signal Y1 :  std_logic_vector(3 downto 0);
   -- timing of Y1: (c0, 0.550000ns)
begin
   with X  select  Y0 <= 
      "0000" when "0000",
      "0001" when "0001",
      "0010" when "0010",
      "0011" when "0011",
      "0100" when "0100",
      "0101" when "0101",
      "0110" when "0110",
      "0111" when "0111",
      "1000" when "1000",
      "1001" when "1001",
      "1010" when "1010",
      "1011" when "1011",
      "1100" when "1100",
      "1101" when "1101",
      "1110" when "1110",
      "1111" when "1111",
      "----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                    LeftShifter11_by_max_20_Freq500_uid4
-- VHDL generated for DummyFPGA @ 500MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca (2008-2011), Florent de Dinechin (2008-2019)
--------------------------------------------------------------------------------
-- Pipeline depth: 1 cycles
-- Clock period (ns): 2
-- Target frequency (MHz): 500
-- Input signals: X S
-- Output signals: R
--  approx. input signal timings: X: (c0, 0.000000ns)S: (c0, 1.090000ns)
--  approx. output signal timings: R: (c1, 1.005385ns)

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity LeftShifter11_by_max_20_Freq500_uid4 is
    port (clk : in std_logic;
          X : in  std_logic_vector(10 downto 0);
          S : in  std_logic_vector(4 downto 0);
          R : out  std_logic_vector(30 downto 0)   );
end entity;

architecture arch of LeftShifter11_by_max_20_Freq500_uid4 is
signal ps, ps_d1 :  std_logic_vector(4 downto 0);
   -- timing of ps: (c0, 1.090000ns)
signal level0 :  std_logic_vector(10 downto 0);
   -- timing of level0: (c0, 0.000000ns)
signal level1, level1_d1 :  std_logic_vector(11 downto 0);
   -- timing of level1: (c0, 1.090000ns)
signal level2 :  std_logic_vector(13 downto 0);
   -- timing of level2: (c1, 0.055385ns)
signal level3 :  std_logic_vector(17 downto 0);
   -- timing of level3: (c1, 0.055385ns)
signal level4 :  std_logic_vector(25 downto 0);
   -- timing of level4: (c1, 1.005385ns)
signal level5 :  std_logic_vector(41 downto 0);
   -- timing of level5: (c1, 1.005385ns)
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            ps_d1 <=  ps;
            level1_d1 <=  level1;
         end if;
      end process;
   ps<= S;
   level0<= X;
   level1<= level0 & (0 downto 0 => '0') when ps(0)= '1' else     (0 downto 0 => '0') & level0;
   level2<= level1_d1 & (1 downto 0 => '0') when ps_d1(1)= '1' else     (1 downto 0 => '0') & level1_d1;
   level3<= level2 & (3 downto 0 => '0') when ps_d1(2)= '1' else     (3 downto 0 => '0') & level2;
   level4<= level3 & (7 downto 0 => '0') when ps_d1(3)= '1' else     (7 downto 0 => '0') & level3;
   level5<= level4 & (15 downto 0 => '0') when ps_d1(4)= '1' else     (15 downto 0 => '0') & level4;
   R <= level5(30 downto 0);
end architecture;

--------------------------------------------------------------------------------
--                         IntAdder_12_Freq500_uid18
-- VHDL generated for DummyFPGA @ 500MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin (2008-2016)
--------------------------------------------------------------------------------
-- Pipeline depth: 2 cycles
-- Clock period (ns): 2
-- Target frequency (MHz): 500
-- Input signals: X Y Cin
-- Output signals: R
--  approx. input signal timings: X: (c1, 1.555385ns)Y: (c1, 1.555385ns)Cin: (c0, 0.000000ns)
--  approx. output signal timings: R: (c2, 0.875385ns)

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntAdder_12_Freq500_uid18 is
    port (clk : in std_logic;
          X : in  std_logic_vector(11 downto 0);
          Y : in  std_logic_vector(11 downto 0);
          Cin : in  std_logic;
          R : out  std_logic_vector(11 downto 0)   );
end entity;

architecture arch of IntAdder_12_Freq500_uid18 is
signal Cin_1, Cin_1_d1, Cin_1_d2 :  std_logic;
   -- timing of Cin_1: (c0, 0.000000ns)
signal X_1, X_1_d1 :  std_logic_vector(12 downto 0);
   -- timing of X_1: (c1, 1.555385ns)
signal Y_1, Y_1_d1 :  std_logic_vector(12 downto 0);
   -- timing of Y_1: (c1, 1.555385ns)
signal S_1 :  std_logic_vector(12 downto 0);
   -- timing of S_1: (c2, 0.875385ns)
signal R_1 :  std_logic_vector(11 downto 0);
   -- timing of R_1: (c2, 0.875385ns)
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            Cin_1_d1 <=  Cin_1;
            Cin_1_d2 <=  Cin_1_d1;
            X_1_d1 <=  X_1;
            Y_1_d1 <=  Y_1;
         end if;
      end process;
   Cin_1 <= Cin;
   X_1 <= '0' & X(11 downto 0);
   Y_1 <= '0' & Y(11 downto 0);
   S_1 <= X_1_d1 + Y_1_d1 + Cin_1_d2;
   R_1 <= S_1(11 downto 0);
   R <= R_1 ;
end architecture;

--------------------------------------------------------------------------------
--                          FixRealKCM_Freq500_uid8
-- VHDL generated for DummyFPGA @ 500MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin (2007-2016)
--------------------------------------------------------------------------------
-- Pipeline depth: 1 cycles
-- Clock period (ns): 2
-- Target frequency (MHz): 500
-- Input signals: X
-- Output signals: R
--  approx. input signal timings: X: (c1, 1.005385ns)
--  approx. output signal timings: R: (c2, 0.875385ns)

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity FixRealKCM_Freq500_uid8 is
    port (clk : in std_logic;
          X : in  std_logic_vector(9 downto 0);
          R : out  std_logic_vector(7 downto 0)   );
end entity;

architecture arch of FixRealKCM_Freq500_uid8 is
   component FixRealKCM_Freq500_uid8_T0_Freq500_uid11 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(11 downto 0)   );
   end component;

   component FixRealKCM_Freq500_uid8_T1_Freq500_uid14 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(6 downto 0)   );
   end component;

   component IntAdder_12_Freq500_uid18 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(11 downto 0);
             Y : in  std_logic_vector(11 downto 0);
             Cin : in  std_logic;
             R : out  std_logic_vector(11 downto 0)   );
   end component;

signal FixRealKCM_Freq500_uid8_A0 :  std_logic_vector(4 downto 0);
   -- timing of FixRealKCM_Freq500_uid8_A0: (c1, 1.005385ns)
signal FixRealKCM_Freq500_uid8_T0 :  std_logic_vector(11 downto 0);
   -- timing of FixRealKCM_Freq500_uid8_T0: (c1, 1.555385ns)
signal FixRealKCM_Freq500_uid8_T0_copy12 :  std_logic_vector(11 downto 0);
   -- timing of FixRealKCM_Freq500_uid8_T0_copy12: (c1, 1.005385ns)
signal bh9_w0_0 :  std_logic;
   -- timing of bh9_w0_0: (c1, 1.555385ns)
signal bh9_w1_0 :  std_logic;
   -- timing of bh9_w1_0: (c1, 1.555385ns)
signal bh9_w2_0 :  std_logic;
   -- timing of bh9_w2_0: (c1, 1.555385ns)
signal bh9_w3_0 :  std_logic;
   -- timing of bh9_w3_0: (c1, 1.555385ns)
signal bh9_w4_0 :  std_logic;
   -- timing of bh9_w4_0: (c1, 1.555385ns)
signal bh9_w5_0 :  std_logic;
   -- timing of bh9_w5_0: (c1, 1.555385ns)
signal bh9_w6_0 :  std_logic;
   -- timing of bh9_w6_0: (c1, 1.555385ns)
signal bh9_w7_0 :  std_logic;
   -- timing of bh9_w7_0: (c1, 1.555385ns)
signal bh9_w8_0 :  std_logic;
   -- timing of bh9_w8_0: (c1, 1.555385ns)
signal bh9_w9_0 :  std_logic;
   -- timing of bh9_w9_0: (c1, 1.555385ns)
signal bh9_w10_0 :  std_logic;
   -- timing of bh9_w10_0: (c1, 1.555385ns)
signal bh9_w11_0 :  std_logic;
   -- timing of bh9_w11_0: (c1, 1.555385ns)
signal FixRealKCM_Freq500_uid8_A1 :  std_logic_vector(4 downto 0);
   -- timing of FixRealKCM_Freq500_uid8_A1: (c1, 1.005385ns)
signal FixRealKCM_Freq500_uid8_T1 :  std_logic_vector(6 downto 0);
   -- timing of FixRealKCM_Freq500_uid8_T1: (c1, 1.555385ns)
signal FixRealKCM_Freq500_uid8_T1_copy15 :  std_logic_vector(6 downto 0);
   -- timing of FixRealKCM_Freq500_uid8_T1_copy15: (c1, 1.005385ns)
signal bh9_w0_1 :  std_logic;
   -- timing of bh9_w0_1: (c1, 1.555385ns)
signal bh9_w1_1 :  std_logic;
   -- timing of bh9_w1_1: (c1, 1.555385ns)
signal bh9_w2_1 :  std_logic;
   -- timing of bh9_w2_1: (c1, 1.555385ns)
signal bh9_w3_1 :  std_logic;
   -- timing of bh9_w3_1: (c1, 1.555385ns)
signal bh9_w4_1 :  std_logic;
   -- timing of bh9_w4_1: (c1, 1.555385ns)
signal bh9_w5_1 :  std_logic;
   -- timing of bh9_w5_1: (c1, 1.555385ns)
signal bh9_w6_1 :  std_logic;
   -- timing of bh9_w6_1: (c1, 1.555385ns)
signal bitheapFinalAdd_bh9_In0 :  std_logic_vector(11 downto 0);
   -- timing of bitheapFinalAdd_bh9_In0: (c1, 1.555385ns)
signal bitheapFinalAdd_bh9_In1 :  std_logic_vector(11 downto 0);
   -- timing of bitheapFinalAdd_bh9_In1: (c1, 1.555385ns)
signal bitheapFinalAdd_bh9_Cin :  std_logic;
   -- timing of bitheapFinalAdd_bh9_Cin: (c0, 0.000000ns)
signal bitheapFinalAdd_bh9_Out :  std_logic_vector(11 downto 0);
   -- timing of bitheapFinalAdd_bh9_Out: (c2, 0.875385ns)
signal bitheapResult_bh9 :  std_logic_vector(11 downto 0);
   -- timing of bitheapResult_bh9: (c2, 0.875385ns)
signal OutRes :  std_logic_vector(11 downto 0);
   -- timing of OutRes: (c2, 0.875385ns)
begin
-- This operator multiplies by 1/log(2)
   FixRealKCM_Freq500_uid8_A0 <= X(9 downto 5);-- input address  m=6  l=2
   FixRealKCM_Freq500_uid8_Table0: FixRealKCM_Freq500_uid8_T0_Freq500_uid11
      port map ( X => FixRealKCM_Freq500_uid8_A0,
                 Y => FixRealKCM_Freq500_uid8_T0_copy12);
   FixRealKCM_Freq500_uid8_T0 <= FixRealKCM_Freq500_uid8_T0_copy12; -- output copy to hold a pipeline register if needed
   bh9_w0_0 <= FixRealKCM_Freq500_uid8_T0(0);
   bh9_w1_0 <= FixRealKCM_Freq500_uid8_T0(1);
   bh9_w2_0 <= FixRealKCM_Freq500_uid8_T0(2);
   bh9_w3_0 <= FixRealKCM_Freq500_uid8_T0(3);
   bh9_w4_0 <= FixRealKCM_Freq500_uid8_T0(4);
   bh9_w5_0 <= FixRealKCM_Freq500_uid8_T0(5);
   bh9_w6_0 <= FixRealKCM_Freq500_uid8_T0(6);
   bh9_w7_0 <= FixRealKCM_Freq500_uid8_T0(7);
   bh9_w8_0 <= FixRealKCM_Freq500_uid8_T0(8);
   bh9_w9_0 <= FixRealKCM_Freq500_uid8_T0(9);
   bh9_w10_0 <= FixRealKCM_Freq500_uid8_T0(10);
   bh9_w11_0 <= FixRealKCM_Freq500_uid8_T0(11);
   FixRealKCM_Freq500_uid8_A1 <= X(4 downto 0);-- input address  m=1  l=-3
   FixRealKCM_Freq500_uid8_Table1: FixRealKCM_Freq500_uid8_T1_Freq500_uid14
      port map ( X => FixRealKCM_Freq500_uid8_A1,
                 Y => FixRealKCM_Freq500_uid8_T1_copy15);
   FixRealKCM_Freq500_uid8_T1 <= FixRealKCM_Freq500_uid8_T1_copy15; -- output copy to hold a pipeline register if needed
   bh9_w0_1 <= FixRealKCM_Freq500_uid8_T1(0);
   bh9_w1_1 <= FixRealKCM_Freq500_uid8_T1(1);
   bh9_w2_1 <= FixRealKCM_Freq500_uid8_T1(2);
   bh9_w3_1 <= FixRealKCM_Freq500_uid8_T1(3);
   bh9_w4_1 <= FixRealKCM_Freq500_uid8_T1(4);
   bh9_w5_1 <= FixRealKCM_Freq500_uid8_T1(5);
   bh9_w6_1 <= FixRealKCM_Freq500_uid8_T1(6);

   -- Adding the constant bits 
      -- All the constant bits are zero, nothing to add


   bitheapFinalAdd_bh9_In0 <= "" & bh9_w11_0 & bh9_w10_0 & bh9_w9_0 & bh9_w8_0 & bh9_w7_0 & bh9_w6_1 & bh9_w5_1 & bh9_w4_1 & bh9_w3_1 & bh9_w2_1 & bh9_w1_1 & bh9_w0_1;
   bitheapFinalAdd_bh9_In1 <= "0" & "0" & "0" & "0" & "0" & bh9_w6_0 & bh9_w5_0 & bh9_w4_0 & bh9_w3_0 & bh9_w2_0 & bh9_w1_0 & bh9_w0_0;
   bitheapFinalAdd_bh9_Cin <= '0';

   bitheapFinalAdd_bh9: IntAdder_12_Freq500_uid18
      port map ( clk  => clk,
                 Cin => bitheapFinalAdd_bh9_Cin,
                 X => bitheapFinalAdd_bh9_In0,
                 Y => bitheapFinalAdd_bh9_In1,
                 R => bitheapFinalAdd_bh9_Out);
   bitheapResult_bh9 <= bitheapFinalAdd_bh9_Out(11 downto 0);
   OutRes <= bitheapResult_bh9(11 downto 0);
   R <= OutRes(11 downto 4);
end architecture;

--------------------------------------------------------------------------------
--                         IntAdder_22_Freq500_uid30
-- VHDL generated for DummyFPGA @ 500MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin (2008-2016)
--------------------------------------------------------------------------------
-- Pipeline depth: 3 cycles
-- Clock period (ns): 2
-- Target frequency (MHz): 500
-- Input signals: X Y Cin
-- Output signals: R
--  approx. input signal timings: X: (c2, 1.425385ns)Y: (c2, 1.425385ns)Cin: (c0, 0.000000ns)
--  approx. output signal timings: R: (c3, 0.835385ns)

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntAdder_22_Freq500_uid30 is
    port (clk : in std_logic;
          X : in  std_logic_vector(21 downto 0);
          Y : in  std_logic_vector(21 downto 0);
          Cin : in  std_logic;
          R : out  std_logic_vector(21 downto 0)   );
end entity;

architecture arch of IntAdder_22_Freq500_uid30 is
signal Rtmp :  std_logic_vector(21 downto 0);
   -- timing of Rtmp: (c3, 0.835385ns)
signal X_d1 :  std_logic_vector(21 downto 0);
   -- timing of X: (c2, 1.425385ns)
signal Y_d1 :  std_logic_vector(21 downto 0);
   -- timing of Y: (c2, 1.425385ns)
signal Cin_d1, Cin_d2, Cin_d3 :  std_logic;
   -- timing of Cin: (c0, 0.000000ns)
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            X_d1 <=  X;
            Y_d1 <=  Y;
            Cin_d1 <=  Cin;
            Cin_d2 <=  Cin_d1;
            Cin_d3 <=  Cin_d2;
         end if;
      end process;
   Rtmp <= X_d1 + Y_d1 + Cin_d3;
   R <= Rtmp;
end architecture;

--------------------------------------------------------------------------------
--                          FixRealKCM_Freq500_uid20
-- VHDL generated for DummyFPGA @ 500MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin (2007-2016)
--------------------------------------------------------------------------------
-- Pipeline depth: 1 cycles
-- Clock period (ns): 2
-- Target frequency (MHz): 500
-- Input signals: X
-- Output signals: R
--  approx. input signal timings: X: (c2, 0.875385ns)
--  approx. output signal timings: R: (c3, 0.835385ns)

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity FixRealKCM_Freq500_uid20 is
    port (clk : in std_logic;
          X : in  std_logic_vector(7 downto 0);
          R : out  std_logic_vector(21 downto 0)   );
end entity;

architecture arch of FixRealKCM_Freq500_uid20 is
   component FixRealKCM_Freq500_uid20_T0_Freq500_uid23 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(21 downto 0)   );
   end component;

   component FixRealKCM_Freq500_uid20_T1_Freq500_uid26 is
      port ( X : in  std_logic_vector(2 downto 0);
             Y : out  std_logic_vector(16 downto 0)   );
   end component;

   component IntAdder_22_Freq500_uid30 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(21 downto 0);
             Y : in  std_logic_vector(21 downto 0);
             Cin : in  std_logic;
             R : out  std_logic_vector(21 downto 0)   );
   end component;

signal FixRealKCM_Freq500_uid20_A0 :  std_logic_vector(4 downto 0);
   -- timing of FixRealKCM_Freq500_uid20_A0: (c2, 0.875385ns)
signal FixRealKCM_Freq500_uid20_T0 :  std_logic_vector(21 downto 0);
   -- timing of FixRealKCM_Freq500_uid20_T0: (c2, 1.425385ns)
signal FixRealKCM_Freq500_uid20_T0_copy24 :  std_logic_vector(21 downto 0);
   -- timing of FixRealKCM_Freq500_uid20_T0_copy24: (c2, 0.875385ns)
signal bh21_w0_0 :  std_logic;
   -- timing of bh21_w0_0: (c2, 1.425385ns)
signal bh21_w1_0 :  std_logic;
   -- timing of bh21_w1_0: (c2, 1.425385ns)
signal bh21_w2_0 :  std_logic;
   -- timing of bh21_w2_0: (c2, 1.425385ns)
signal bh21_w3_0 :  std_logic;
   -- timing of bh21_w3_0: (c2, 1.425385ns)
signal bh21_w4_0 :  std_logic;
   -- timing of bh21_w4_0: (c2, 1.425385ns)
signal bh21_w5_0 :  std_logic;
   -- timing of bh21_w5_0: (c2, 1.425385ns)
signal bh21_w6_0 :  std_logic;
   -- timing of bh21_w6_0: (c2, 1.425385ns)
signal bh21_w7_0 :  std_logic;
   -- timing of bh21_w7_0: (c2, 1.425385ns)
signal bh21_w8_0 :  std_logic;
   -- timing of bh21_w8_0: (c2, 1.425385ns)
signal bh21_w9_0 :  std_logic;
   -- timing of bh21_w9_0: (c2, 1.425385ns)
signal bh21_w10_0 :  std_logic;
   -- timing of bh21_w10_0: (c2, 1.425385ns)
signal bh21_w11_0 :  std_logic;
   -- timing of bh21_w11_0: (c2, 1.425385ns)
signal bh21_w12_0 :  std_logic;
   -- timing of bh21_w12_0: (c2, 1.425385ns)
signal bh21_w13_0 :  std_logic;
   -- timing of bh21_w13_0: (c2, 1.425385ns)
signal bh21_w14_0 :  std_logic;
   -- timing of bh21_w14_0: (c2, 1.425385ns)
signal bh21_w15_0 :  std_logic;
   -- timing of bh21_w15_0: (c2, 1.425385ns)
signal bh21_w16_0 :  std_logic;
   -- timing of bh21_w16_0: (c2, 1.425385ns)
signal bh21_w17_0 :  std_logic;
   -- timing of bh21_w17_0: (c2, 1.425385ns)
signal bh21_w18_0 :  std_logic;
   -- timing of bh21_w18_0: (c2, 1.425385ns)
signal bh21_w19_0 :  std_logic;
   -- timing of bh21_w19_0: (c2, 1.425385ns)
signal bh21_w20_0 :  std_logic;
   -- timing of bh21_w20_0: (c2, 1.425385ns)
signal bh21_w21_0 :  std_logic;
   -- timing of bh21_w21_0: (c2, 1.425385ns)
signal FixRealKCM_Freq500_uid20_A1 :  std_logic_vector(2 downto 0);
   -- timing of FixRealKCM_Freq500_uid20_A1: (c2, 0.875385ns)
signal FixRealKCM_Freq500_uid20_T1 :  std_logic_vector(16 downto 0);
   -- timing of FixRealKCM_Freq500_uid20_T1: (c2, 1.425385ns)
signal FixRealKCM_Freq500_uid20_T1_copy27 :  std_logic_vector(16 downto 0);
   -- timing of FixRealKCM_Freq500_uid20_T1_copy27: (c2, 0.875385ns)
signal bh21_w0_1 :  std_logic;
   -- timing of bh21_w0_1: (c2, 1.425385ns)
signal bh21_w1_1 :  std_logic;
   -- timing of bh21_w1_1: (c2, 1.425385ns)
signal bh21_w2_1 :  std_logic;
   -- timing of bh21_w2_1: (c2, 1.425385ns)
signal bh21_w3_1 :  std_logic;
   -- timing of bh21_w3_1: (c2, 1.425385ns)
signal bh21_w4_1 :  std_logic;
   -- timing of bh21_w4_1: (c2, 1.425385ns)
signal bh21_w5_1 :  std_logic;
   -- timing of bh21_w5_1: (c2, 1.425385ns)
signal bh21_w6_1 :  std_logic;
   -- timing of bh21_w6_1: (c2, 1.425385ns)
signal bh21_w7_1 :  std_logic;
   -- timing of bh21_w7_1: (c2, 1.425385ns)
signal bh21_w8_1 :  std_logic;
   -- timing of bh21_w8_1: (c2, 1.425385ns)
signal bh21_w9_1 :  std_logic;
   -- timing of bh21_w9_1: (c2, 1.425385ns)
signal bh21_w10_1 :  std_logic;
   -- timing of bh21_w10_1: (c2, 1.425385ns)
signal bh21_w11_1 :  std_logic;
   -- timing of bh21_w11_1: (c2, 1.425385ns)
signal bh21_w12_1 :  std_logic;
   -- timing of bh21_w12_1: (c2, 1.425385ns)
signal bh21_w13_1 :  std_logic;
   -- timing of bh21_w13_1: (c2, 1.425385ns)
signal bh21_w14_1 :  std_logic;
   -- timing of bh21_w14_1: (c2, 1.425385ns)
signal bh21_w15_1 :  std_logic;
   -- timing of bh21_w15_1: (c2, 1.425385ns)
signal bh21_w16_1 :  std_logic;
   -- timing of bh21_w16_1: (c2, 1.425385ns)
signal bitheapFinalAdd_bh21_In0 :  std_logic_vector(21 downto 0);
   -- timing of bitheapFinalAdd_bh21_In0: (c2, 1.425385ns)
signal bitheapFinalAdd_bh21_In1 :  std_logic_vector(21 downto 0);
   -- timing of bitheapFinalAdd_bh21_In1: (c2, 1.425385ns)
signal bitheapFinalAdd_bh21_Cin :  std_logic;
   -- timing of bitheapFinalAdd_bh21_Cin: (c0, 0.000000ns)
signal bitheapFinalAdd_bh21_Out :  std_logic_vector(21 downto 0);
   -- timing of bitheapFinalAdd_bh21_Out: (c3, 0.835385ns)
signal bitheapResult_bh21 :  std_logic_vector(21 downto 0);
   -- timing of bitheapResult_bh21: (c3, 0.835385ns)
signal OutRes :  std_logic_vector(21 downto 0);
   -- timing of OutRes: (c3, 0.835385ns)
begin
-- This operator multiplies by log(2)
   FixRealKCM_Freq500_uid20_A0 <= X(7 downto 3);-- input address  m=7  l=3
   FixRealKCM_Freq500_uid20_Table0: FixRealKCM_Freq500_uid20_T0_Freq500_uid23
      port map ( X => FixRealKCM_Freq500_uid20_A0,
                 Y => FixRealKCM_Freq500_uid20_T0_copy24);
   FixRealKCM_Freq500_uid20_T0 <= FixRealKCM_Freq500_uid20_T0_copy24; -- output copy to hold a pipeline register if needed
   bh21_w0_0 <= FixRealKCM_Freq500_uid20_T0(0);
   bh21_w1_0 <= FixRealKCM_Freq500_uid20_T0(1);
   bh21_w2_0 <= FixRealKCM_Freq500_uid20_T0(2);
   bh21_w3_0 <= FixRealKCM_Freq500_uid20_T0(3);
   bh21_w4_0 <= FixRealKCM_Freq500_uid20_T0(4);
   bh21_w5_0 <= FixRealKCM_Freq500_uid20_T0(5);
   bh21_w6_0 <= FixRealKCM_Freq500_uid20_T0(6);
   bh21_w7_0 <= FixRealKCM_Freq500_uid20_T0(7);
   bh21_w8_0 <= FixRealKCM_Freq500_uid20_T0(8);
   bh21_w9_0 <= FixRealKCM_Freq500_uid20_T0(9);
   bh21_w10_0 <= FixRealKCM_Freq500_uid20_T0(10);
   bh21_w11_0 <= FixRealKCM_Freq500_uid20_T0(11);
   bh21_w12_0 <= FixRealKCM_Freq500_uid20_T0(12);
   bh21_w13_0 <= FixRealKCM_Freq500_uid20_T0(13);
   bh21_w14_0 <= FixRealKCM_Freq500_uid20_T0(14);
   bh21_w15_0 <= FixRealKCM_Freq500_uid20_T0(15);
   bh21_w16_0 <= FixRealKCM_Freq500_uid20_T0(16);
   bh21_w17_0 <= FixRealKCM_Freq500_uid20_T0(17);
   bh21_w18_0 <= FixRealKCM_Freq500_uid20_T0(18);
   bh21_w19_0 <= FixRealKCM_Freq500_uid20_T0(19);
   bh21_w20_0 <= FixRealKCM_Freq500_uid20_T0(20);
   bh21_w21_0 <= FixRealKCM_Freq500_uid20_T0(21);
   FixRealKCM_Freq500_uid20_A1 <= X(2 downto 0);-- input address  m=2  l=0
   FixRealKCM_Freq500_uid20_Table1: FixRealKCM_Freq500_uid20_T1_Freq500_uid26
      port map ( X => FixRealKCM_Freq500_uid20_A1,
                 Y => FixRealKCM_Freq500_uid20_T1_copy27);
   FixRealKCM_Freq500_uid20_T1 <= FixRealKCM_Freq500_uid20_T1_copy27; -- output copy to hold a pipeline register if needed
   bh21_w0_1 <= FixRealKCM_Freq500_uid20_T1(0);
   bh21_w1_1 <= FixRealKCM_Freq500_uid20_T1(1);
   bh21_w2_1 <= FixRealKCM_Freq500_uid20_T1(2);
   bh21_w3_1 <= FixRealKCM_Freq500_uid20_T1(3);
   bh21_w4_1 <= FixRealKCM_Freq500_uid20_T1(4);
   bh21_w5_1 <= FixRealKCM_Freq500_uid20_T1(5);
   bh21_w6_1 <= FixRealKCM_Freq500_uid20_T1(6);
   bh21_w7_1 <= FixRealKCM_Freq500_uid20_T1(7);
   bh21_w8_1 <= FixRealKCM_Freq500_uid20_T1(8);
   bh21_w9_1 <= FixRealKCM_Freq500_uid20_T1(9);
   bh21_w10_1 <= FixRealKCM_Freq500_uid20_T1(10);
   bh21_w11_1 <= FixRealKCM_Freq500_uid20_T1(11);
   bh21_w12_1 <= FixRealKCM_Freq500_uid20_T1(12);
   bh21_w13_1 <= FixRealKCM_Freq500_uid20_T1(13);
   bh21_w14_1 <= FixRealKCM_Freq500_uid20_T1(14);
   bh21_w15_1 <= FixRealKCM_Freq500_uid20_T1(15);
   bh21_w16_1 <= FixRealKCM_Freq500_uid20_T1(16);

   -- Adding the constant bits 
      -- All the constant bits are zero, nothing to add


   bitheapFinalAdd_bh21_In0 <= "" & bh21_w21_0 & bh21_w20_0 & bh21_w19_0 & bh21_w18_0 & bh21_w17_0 & bh21_w16_0 & bh21_w15_0 & bh21_w14_0 & bh21_w13_0 & bh21_w12_0 & bh21_w11_0 & bh21_w10_0 & bh21_w9_0 & bh21_w8_0 & bh21_w7_0 & bh21_w6_0 & bh21_w5_0 & bh21_w4_0 & bh21_w3_0 & bh21_w2_0 & bh21_w1_0 & bh21_w0_0;
   bitheapFinalAdd_bh21_In1 <= "0" & "0" & "0" & "0" & "0" & bh21_w16_1 & bh21_w15_1 & bh21_w14_1 & bh21_w13_1 & bh21_w12_1 & bh21_w11_1 & bh21_w10_1 & bh21_w9_1 & bh21_w8_1 & bh21_w7_1 & bh21_w6_1 & bh21_w5_1 & bh21_w4_1 & bh21_w3_1 & bh21_w2_1 & bh21_w1_1 & bh21_w0_1;
   bitheapFinalAdd_bh21_Cin <= '0';

   bitheapFinalAdd_bh21: IntAdder_22_Freq500_uid30
      port map ( clk  => clk,
                 Cin => bitheapFinalAdd_bh21_Cin,
                 X => bitheapFinalAdd_bh21_In0,
                 Y => bitheapFinalAdd_bh21_In1,
                 R => bitheapFinalAdd_bh21_Out);
   bitheapResult_bh21 <= bitheapFinalAdd_bh21_Out(21 downto 0);
   OutRes <= bitheapResult_bh21(21 downto 0);
   R <= OutRes(21 downto 0);
end architecture;

--------------------------------------------------------------------------------
--                         IntAdder_14_Freq500_uid33
-- VHDL generated for DummyFPGA @ 500MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin (2008-2016)
--------------------------------------------------------------------------------
-- Pipeline depth: 4 cycles
-- Clock period (ns): 2
-- Target frequency (MHz): 500
-- Input signals: X Y Cin
-- Output signals: R
--  approx. input signal timings: X: (c1, 1.555385ns)Y: (c3, 0.835385ns)Cin: (c0, 0.000000ns)
--  approx. output signal timings: R: (c4, 0.175385ns)

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntAdder_14_Freq500_uid33 is
    port (clk : in std_logic;
          X : in  std_logic_vector(13 downto 0);
          Y : in  std_logic_vector(13 downto 0);
          Cin : in  std_logic;
          R : out  std_logic_vector(13 downto 0)   );
end entity;

architecture arch of IntAdder_14_Freq500_uid33 is
signal Cin_1, Cin_1_d1, Cin_1_d2, Cin_1_d3, Cin_1_d4 :  std_logic;
   -- timing of Cin_1: (c0, 0.000000ns)
signal X_1, X_1_d1, X_1_d2, X_1_d3 :  std_logic_vector(14 downto 0);
   -- timing of X_1: (c1, 1.555385ns)
signal Y_1, Y_1_d1 :  std_logic_vector(14 downto 0);
   -- timing of Y_1: (c3, 0.835385ns)
signal S_1 :  std_logic_vector(14 downto 0);
   -- timing of S_1: (c4, 0.175385ns)
signal R_1 :  std_logic_vector(13 downto 0);
   -- timing of R_1: (c4, 0.175385ns)
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            Cin_1_d1 <=  Cin_1;
            Cin_1_d2 <=  Cin_1_d1;
            Cin_1_d3 <=  Cin_1_d2;
            Cin_1_d4 <=  Cin_1_d3;
            X_1_d1 <=  X_1;
            X_1_d2 <=  X_1_d1;
            X_1_d3 <=  X_1_d2;
            Y_1_d1 <=  Y_1;
         end if;
      end process;
   Cin_1 <= Cin;
   X_1 <= '0' & X(13 downto 0);
   Y_1 <= '0' & Y(13 downto 0);
   S_1 <= X_1_d3 + Y_1_d1 + Cin_1_d4;
   R_1 <= S_1(13 downto 0);
   R <= R_1 ;
end architecture;

--------------------------------------------------------------------------------
--                          IntAdder_5_Freq500_uid43
-- VHDL generated for DummyFPGA @ 500MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin (2008-2016)
--------------------------------------------------------------------------------
-- Pipeline depth: 4 cycles
-- Clock period (ns): 2
-- Target frequency (MHz): 500
-- Input signals: X Y Cin
-- Output signals: R
--  approx. input signal timings: X: (c4, 0.725385ns)Y: (c0, 0.000000ns)Cin: (c0, 0.000000ns)
--  approx. output signal timings: R: (c4, 1.765385ns)

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntAdder_5_Freq500_uid43 is
    port (clk : in std_logic;
          X : in  std_logic_vector(4 downto 0);
          Y : in  std_logic_vector(4 downto 0);
          Cin : in  std_logic;
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntAdder_5_Freq500_uid43 is
signal Rtmp :  std_logic_vector(4 downto 0);
   -- timing of Rtmp: (c4, 1.765385ns)
signal Y_d1, Y_d2, Y_d3, Y_d4 :  std_logic_vector(4 downto 0);
   -- timing of Y: (c0, 0.000000ns)
signal Cin_d1, Cin_d2, Cin_d3, Cin_d4 :  std_logic;
   -- timing of Cin: (c0, 0.000000ns)
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            Y_d1 <=  Y;
            Y_d2 <=  Y_d1;
            Y_d3 <=  Y_d2;
            Y_d4 <=  Y_d3;
            Cin_d1 <=  Cin;
            Cin_d2 <=  Cin_d1;
            Cin_d3 <=  Cin_d2;
            Cin_d4 <=  Cin_d3;
         end if;
      end process;
   Rtmp <= X + Y_d4 + Cin_d4;
   R <= Rtmp;
end architecture;

--------------------------------------------------------------------------------
--                     IntMultiplier_4x5_6_Freq500_uid45
-- VHDL generated for DummyFPGA @ 500MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Martin Kumm, Florent de Dinechin, Andreas Böttcher, Kinga Illyes, Bogdan Popa, Bogdan Pasca, 2012-
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 2
-- Target frequency (MHz): 500
-- Input signals: X Y
-- Output signals: R
--  approx. input signal timings: X: (c4, 1.765385ns)Y: (c4, 0.725385ns)
--  approx. output signal timings: R: (c4, 1.765385ns)

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity IntMultiplier_4x5_6_Freq500_uid45 is
    port (clk : in std_logic;
          X : in  std_logic_vector(3 downto 0);
          Y : in  std_logic_vector(4 downto 0);
          R : out  std_logic_vector(5 downto 0)   );
end entity;

architecture arch of IntMultiplier_4x5_6_Freq500_uid45 is
signal XX_m46 :  std_logic_vector(3 downto 0);
   -- timing of XX_m46: (c4, 1.765385ns)
signal YY_m46 :  std_logic_vector(4 downto 0);
   -- timing of YY_m46: (c4, 0.725385ns)
signal XX :  unsigned(-1+4 downto 0);
   -- timing of XX: (c4, 1.765385ns)
signal YY :  unsigned(-1+5 downto 0);
   -- timing of YY: (c4, 0.725385ns)
signal RR :  unsigned(-1+9 downto 0);
   -- timing of RR: (c4, 1.765385ns)
begin
   XX_m46 <= X ;
   YY_m46 <= Y ;
   XX <= unsigned(X);
   YY <= unsigned(Y);
   RR <= XX*YY;
   R <= std_logic_vector(RR(8 downto 3));
end architecture;

--------------------------------------------------------------------------------
--                         IntAdder_15_Freq500_uid49
-- VHDL generated for DummyFPGA @ 500MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin (2008-2016)
--------------------------------------------------------------------------------
-- Pipeline depth: 5 cycles
-- Clock period (ns): 2
-- Target frequency (MHz): 500
-- Input signals: X Y Cin
-- Output signals: R
--  approx. input signal timings: X: (c4, 0.725385ns)Y: (c4, 1.765385ns)Cin: (c0, 0.000000ns)
--  approx. output signal timings: R: (c5, 1.105385ns)

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntAdder_15_Freq500_uid49 is
    port (clk : in std_logic;
          X : in  std_logic_vector(14 downto 0);
          Y : in  std_logic_vector(14 downto 0);
          Cin : in  std_logic;
          R : out  std_logic_vector(14 downto 0)   );
end entity;

architecture arch of IntAdder_15_Freq500_uid49 is
signal Rtmp :  std_logic_vector(14 downto 0);
   -- timing of Rtmp: (c5, 1.105385ns)
signal X_d1 :  std_logic_vector(14 downto 0);
   -- timing of X: (c4, 0.725385ns)
signal Y_d1 :  std_logic_vector(14 downto 0);
   -- timing of Y: (c4, 1.765385ns)
signal Cin_d1, Cin_d2, Cin_d3, Cin_d4, Cin_d5 :  std_logic;
   -- timing of Cin: (c0, 0.000000ns)
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            X_d1 <=  X;
            Y_d1 <=  Y;
            Cin_d1 <=  Cin;
            Cin_d2 <=  Cin_d1;
            Cin_d3 <=  Cin_d2;
            Cin_d4 <=  Cin_d3;
            Cin_d5 <=  Cin_d4;
         end if;
      end process;
   Rtmp <= X_d1 + Y_d1 + Cin_d5;
   R <= Rtmp;
end architecture;

--------------------------------------------------------------------------------
--                           Exp_8_10_Freq500_uid6
-- VHDL generated for DummyFPGA @ 500MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: F. de Dinechin, Bogdan Pasca, Orégane Desrentes (2008-2025)
--------------------------------------------------------------------------------
-- Pipeline depth: 5 cycles
-- Clock period (ns): 2
-- Target frequency (MHz): 500
-- Input signals: ufixX_i XSign
-- Output signals: expY K
--  approx. input signal timings: ufixX_i: (c1, 1.005385ns)XSign: (c0, 0.000000ns)
--  approx. output signal timings: expY: (c5, 1.105385ns)K: (c3, 0.155385ns)

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity Exp_8_10_Freq500_uid6 is
    port (clk : in std_logic;
          ufixX_i : in  std_logic_vector(20 downto 0);
          XSign : in  std_logic;
          expY : out  std_logic_vector(14 downto 0);
          K : out  std_logic_vector(8 downto 0)   );
end entity;

architecture arch of Exp_8_10_Freq500_uid6 is
   component FixRealKCM_Freq500_uid8 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(9 downto 0);
             R : out  std_logic_vector(7 downto 0)   );
   end component;

   component FixRealKCM_Freq500_uid20 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(7 downto 0);
             R : out  std_logic_vector(21 downto 0)   );
   end component;

   component IntAdder_14_Freq500_uid33 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(13 downto 0);
             Y : in  std_logic_vector(13 downto 0);
             Cin : in  std_logic;
             R : out  std_logic_vector(13 downto 0)   );
   end component;

   component FixFunctionByTable_Freq500_uid35 is
      port ( X : in  std_logic_vector(9 downto 0);
             Y : out  std_logic_vector(14 downto 0)   );
   end component;

   component FixFunctionByTable_Freq500_uid38 is
      port ( X : in  std_logic_vector(3 downto 0);
             Y : out  std_logic_vector(3 downto 0)   );
   end component;

   component IntAdder_5_Freq500_uid43 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(4 downto 0);
             Y : in  std_logic_vector(4 downto 0);
             Cin : in  std_logic;
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplier_4x5_6_Freq500_uid45 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(3 downto 0);
             Y : in  std_logic_vector(4 downto 0);
             R : out  std_logic_vector(5 downto 0)   );
   end component;

   component IntAdder_15_Freq500_uid49 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(14 downto 0);
             Y : in  std_logic_vector(14 downto 0);
             Cin : in  std_logic;
             R : out  std_logic_vector(14 downto 0)   );
   end component;

signal ufixX :  unsigned(6+14 downto 0);
   -- timing of ufixX: (c1, 1.005385ns)
signal xMulIn :  unsigned(6+3 downto 0);
   -- timing of xMulIn: (c1, 1.005385ns)
signal absK, absK_d1 :  std_logic_vector(7 downto 0);
   -- timing of absK: (c2, 0.875385ns)
signal minusAbsK :  std_logic_vector(8 downto 0);
   -- timing of minusAbsK: (c3, 0.155385ns)
signal absKLog2 :  std_logic_vector(21 downto 0);
   -- timing of absKLog2: (c3, 0.835385ns)
signal subOp1 :  std_logic_vector(13 downto 0);
   -- timing of subOp1: (c1, 1.555385ns)
signal subOp2 :  std_logic_vector(13 downto 0);
   -- timing of subOp2: (c3, 0.835385ns)
signal Y :  std_logic_vector(13 downto 0);
   -- timing of Y: (c4, 0.175385ns)
signal A :  std_logic_vector(9 downto 0);
   -- timing of A: (c4, 0.175385ns)
signal Z :  std_logic_vector(3 downto 0);
   -- timing of Z: (c4, 0.175385ns)
signal expA :  std_logic_vector(14 downto 0);
   -- timing of expA: (c4, 0.725385ns)
signal expA_copy36 :  std_logic_vector(14 downto 0);
   -- timing of expA_copy36: (c4, 0.175385ns)
signal expZm1_p :  std_logic_vector(3 downto 0);
   -- timing of expZm1_p: (c4, 0.725385ns)
signal expZm1_p_copy39 :  std_logic_vector(3 downto 0);
   -- timing of expZm1_p_copy39: (c4, 0.175385ns)
signal expZm1 :  std_logic_vector(4 downto 0);
   -- timing of expZm1: (c4, 0.725385ns)
signal expA_T :  std_logic_vector(4 downto 0);
   -- timing of expA_T: (c4, 0.725385ns)
signal expArounded0 :  std_logic_vector(4 downto 0);
   -- timing of expArounded0: (c4, 1.765385ns)
signal expArounded :  std_logic_vector(3 downto 0);
   -- timing of expArounded: (c4, 1.765385ns)
signal lowerProduct :  std_logic_vector(5 downto 0);
   -- timing of lowerProduct: (c4, 1.765385ns)
signal extendedLowerProduct :  std_logic_vector(14 downto 0);
   -- timing of extendedLowerProduct: (c4, 1.765385ns)
signal XSign_d1, XSign_d2, XSign_d3 :  std_logic;
   -- timing of XSign: (c0, 0.000000ns)
constant g: positive := 4;
constant wE: positive := 8;
constant wF: positive := 10;
constant wFIn: positive := 10;
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            absK_d1 <=  absK;
            XSign_d1 <=  XSign;
            XSign_d2 <=  XSign_d1;
            XSign_d3 <=  XSign_d2;
         end if;
      end process;
ufixX <= unsigned(ufixX_i);
   xMulIn <= ufixX(20 downto 11); -- fix resize from (6, -14) to (6, -3)
   MulInvLog2: FixRealKCM_Freq500_uid8
      port map ( clk  => clk,
                 X => std_logic_vector(xMulIn),
                 R => absK);
   minusAbsK <= (8 downto 0 => '0') - ('0' & absK_d1);
   K <= minusAbsK when  XSign_d3='1'   else ('0' & absK_d1);
   MulLog2: FixRealKCM_Freq500_uid20
      port map ( clk  => clk,
                 X => absK,
                 R => absKLog2);
   subOp1 <= std_logic_vector(ufixX(13 downto 0)) when XSign_d1='0' else not (std_logic_vector(ufixX(13 downto 0)));
   subOp2 <= absKLog2(13 downto 0) when XSign_d3='1' else not (absKLog2(13 downto 0));
   theYAdder: IntAdder_14_Freq500_uid33
      port map ( clk  => clk,
                 Cin => '1',
                 X => subOp1,
                 Y => subOp2,
                 R => Y);
   -- Now compute the exp of this fixed-point value
   A <= Y(13 downto 4);
   Z <= Y(3 downto 0);
   ExpATable: FixFunctionByTable_Freq500_uid35
      port map ( X => A,
                 Y => expA_copy36);
   expA <= expA_copy36; -- output copy to hold a pipeline register if needed
   ExpZm1Table: FixFunctionByTable_Freq500_uid38
      port map ( X => Z,
                 Y => expZm1_p_copy39);
   expZm1_p <= expZm1_p_copy39; -- output copy to hold a pipeline register if needed
expZm1 <= "0" & expZm1_p;
   -- Rounding expA to the same accuracy as expZm1
   --   (truncation would not be accurate enough and require one more guard bit)
   expA_T <= expA(14 downto 10);
   Adder_expArounded0: IntAdder_5_Freq500_uid43
      port map ( clk  => clk,
                 Cin => '1',
                 X => expA_T,
                 Y => "00000",
                 R => expArounded0);
   expArounded <= expArounded0(4 downto 1);
   TheLowerProduct: IntMultiplier_4x5_6_Freq500_uid45
      port map ( clk  => clk,
                 X => expArounded,
                 Y => expZm1,
                 R => lowerProduct);
   extendedLowerProduct <= ((14 downto 6 => '0') & lowerProduct(5 downto 0));
   -- Final addition -- the product MSB bit weight is -k+2 = -8
   TheFinalAdder: IntAdder_15_Freq500_uid49
      port map ( clk  => clk,
                 Cin => '0',
                 X => expA,
                 Y => extendedLowerProduct,
                 R => expY);
end architecture;

--------------------------------------------------------------------------------
--                         IntAdder_20_Freq500_uid52
-- VHDL generated for DummyFPGA @ 500MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin (2008-2016)
--------------------------------------------------------------------------------
-- Pipeline depth: 6 cycles
-- Clock period (ns): 2
-- Target frequency (MHz): 500
-- Input signals: X Y Cin
-- Output signals: R
--  approx. input signal timings: X: (c5, 1.655385ns)Y: (c5, 1.105385ns)Cin: (c0, 0.000000ns)
--  approx. output signal timings: R: (c6, 1.055385ns)

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntAdder_20_Freq500_uid52 is
    port (clk : in std_logic;
          X : in  std_logic_vector(19 downto 0);
          Y : in  std_logic_vector(19 downto 0);
          Cin : in  std_logic;
          R : out  std_logic_vector(19 downto 0)   );
end entity;

architecture arch of IntAdder_20_Freq500_uid52 is
signal Cin_1, Cin_1_d1, Cin_1_d2, Cin_1_d3, Cin_1_d4, Cin_1_d5, Cin_1_d6 :  std_logic;
   -- timing of Cin_1: (c0, 0.000000ns)
signal X_1, X_1_d1 :  std_logic_vector(20 downto 0);
   -- timing of X_1: (c5, 1.655385ns)
signal Y_1, Y_1_d1 :  std_logic_vector(20 downto 0);
   -- timing of Y_1: (c5, 1.105385ns)
signal S_1 :  std_logic_vector(20 downto 0);
   -- timing of S_1: (c6, 1.055385ns)
signal R_1 :  std_logic_vector(19 downto 0);
   -- timing of R_1: (c6, 1.055385ns)
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            Cin_1_d1 <=  Cin_1;
            Cin_1_d2 <=  Cin_1_d1;
            Cin_1_d3 <=  Cin_1_d2;
            Cin_1_d4 <=  Cin_1_d3;
            Cin_1_d5 <=  Cin_1_d4;
            Cin_1_d6 <=  Cin_1_d5;
            X_1_d1 <=  X_1;
            Y_1_d1 <=  Y_1;
         end if;
      end process;
   Cin_1 <= Cin;
   X_1 <= '0' & X(19 downto 0);
   Y_1 <= '0' & Y(19 downto 0);
   S_1 <= X_1_d1 + Y_1_d1 + Cin_1_d6;
   R_1 <= S_1(19 downto 0);
   R <= R_1 ;
end architecture;

--------------------------------------------------------------------------------
--                                 top_module
--                         (FPExp_8_10_Freq500_uid2)
-- VHDL generated for DummyFPGA @ 500MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: F. de Dinechin, Bogdan Pasca, Orégane Desrentes (2008-2025)
--------------------------------------------------------------------------------
-- Pipeline depth: 6 cycles
-- Clock period (ns): 2
-- Target frequency (MHz): 500
-- Input signals: X
-- Output signals: R
--  approx. input signal timings: X: (c0, 0.000000ns)
--  approx. output signal timings: R: (c6, 1.605385ns)

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity top_module is
    port (clk : in std_logic;
          X : in  std_logic_vector(8+10+2 downto 0);
          R : out  std_logic_vector(8+10+2 downto 0)   );
end entity;

architecture arch of top_module is
   component LeftShifter11_by_max_20_Freq500_uid4 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(10 downto 0);
             S : in  std_logic_vector(4 downto 0);
             R : out  std_logic_vector(30 downto 0)   );
   end component;

   component Exp_8_10_Freq500_uid6 is
      port ( clk : in std_logic;
             ufixX_i : in  std_logic_vector(20 downto 0);
             XSign : in  std_logic;
             expY : out  std_logic_vector(14 downto 0);
             K : out  std_logic_vector(8 downto 0)   );
   end component;

   component IntAdder_20_Freq500_uid52 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(19 downto 0);
             Y : in  std_logic_vector(19 downto 0);
             Cin : in  std_logic;
             R : out  std_logic_vector(19 downto 0)   );
   end component;

signal Xexn, Xexn_d1, Xexn_d2, Xexn_d3, Xexn_d4, Xexn_d5, Xexn_d6 :  std_logic_vector(1 downto 0);
   -- timing of Xexn: (c0, 0.000000ns)
signal XSign, XSign_d1, XSign_d2, XSign_d3, XSign_d4, XSign_d5, XSign_d6 :  std_logic;
   -- timing of XSign: (c0, 0.000000ns)
signal XexpField :  std_logic_vector(7 downto 0);
   -- timing of XexpField: (c0, 0.000000ns)
signal Xfrac :  unsigned(-1+10 downto 0);
   -- timing of Xfrac: (c0, 0.000000ns)
signal e0 :  std_logic_vector(9 downto 0);
   -- timing of e0: (c0, 0.000000ns)
signal shiftVal, shiftVal_d1 :  std_logic_vector(9 downto 0);
   -- timing of shiftVal: (c0, 1.090000ns)
signal resultWillBeOne, resultWillBeOne_d1 :  std_logic;
   -- timing of resultWillBeOne: (c0, 1.090000ns)
signal mXu :  unsigned(0+10 downto 0);
   -- timing of mXu: (c0, 0.000000ns)
signal maxShift, maxShift_d1 :  std_logic_vector(8 downto 0);
   -- timing of maxShift: (c0, 0.000000ns)
signal overflow0 :  std_logic;
   -- timing of overflow0: (c1, 0.370000ns)
signal shiftValIn :  std_logic_vector(4 downto 0);
   -- timing of shiftValIn: (c0, 1.090000ns)
signal fixX0 :  std_logic_vector(30 downto 0);
   -- timing of fixX0: (c1, 1.005385ns)
signal ufixX :  unsigned(6+14 downto 0);
   -- timing of ufixX: (c1, 1.005385ns)
signal expY :  std_logic_vector(14 downto 0);
   -- timing of expY: (c5, 1.105385ns)
signal K, K_d1, K_d2 :  std_logic_vector(8 downto 0);
   -- timing of K: (c3, 0.155385ns)
signal needNoNorm :  std_logic;
   -- timing of needNoNorm: (c5, 1.105385ns)
signal preRoundBiasSig :  std_logic_vector(19 downto 0);
   -- timing of preRoundBiasSig: (c5, 1.655385ns)
signal roundBit :  std_logic;
   -- timing of roundBit: (c5, 1.105385ns)
signal roundNormAddend :  std_logic_vector(19 downto 0);
   -- timing of roundNormAddend: (c5, 1.105385ns)
signal roundedExpSigRes :  std_logic_vector(19 downto 0);
   -- timing of roundedExpSigRes: (c6, 1.055385ns)
signal roundedExpSig :  std_logic_vector(19 downto 0);
   -- timing of roundedExpSig: (c6, 1.605385ns)
signal ofl1, ofl1_d1, ofl1_d2, ofl1_d3, ofl1_d4, ofl1_d5 :  std_logic;
   -- timing of ofl1: (c1, 0.920000ns)
signal ofl2 :  std_logic;
   -- timing of ofl2: (c6, 1.605385ns)
signal ofl3, ofl3_d1, ofl3_d2, ofl3_d3, ofl3_d4, ofl3_d5, ofl3_d6 :  std_logic;
   -- timing of ofl3: (c0, 0.000000ns)
signal ofl :  std_logic;
   -- timing of ofl: (c6, 1.605385ns)
signal ufl1 :  std_logic;
   -- timing of ufl1: (c6, 1.605385ns)
signal ufl2, ufl2_d1, ufl2_d2, ufl2_d3, ufl2_d4, ufl2_d5, ufl2_d6 :  std_logic;
   -- timing of ufl2: (c0, 0.000000ns)
signal ufl3, ufl3_d1, ufl3_d2, ufl3_d3, ufl3_d4, ufl3_d5 :  std_logic;
   -- timing of ufl3: (c1, 0.370000ns)
signal ufl :  std_logic;
   -- timing of ufl: (c6, 1.605385ns)
signal Rexn :  std_logic_vector(1 downto 0);
   -- timing of Rexn: (c6, 1.605385ns)
constant g: positive := 4;
constant wE: positive := 8;
constant wF: positive := 10;
constant wFIn: positive := 10;
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            Xexn_d1 <=  Xexn;
            Xexn_d2 <=  Xexn_d1;
            Xexn_d3 <=  Xexn_d2;
            Xexn_d4 <=  Xexn_d3;
            Xexn_d5 <=  Xexn_d4;
            Xexn_d6 <=  Xexn_d5;
            XSign_d1 <=  XSign;
            XSign_d2 <=  XSign_d1;
            XSign_d3 <=  XSign_d2;
            XSign_d4 <=  XSign_d3;
            XSign_d5 <=  XSign_d4;
            XSign_d6 <=  XSign_d5;
            shiftVal_d1 <=  shiftVal;
            resultWillBeOne_d1 <=  resultWillBeOne;
            maxShift_d1 <=  maxShift;
            K_d1 <=  K;
            K_d2 <=  K_d1;
            ofl1_d1 <=  ofl1;
            ofl1_d2 <=  ofl1_d1;
            ofl1_d3 <=  ofl1_d2;
            ofl1_d4 <=  ofl1_d3;
            ofl1_d5 <=  ofl1_d4;
            ofl3_d1 <=  ofl3;
            ofl3_d2 <=  ofl3_d1;
            ofl3_d3 <=  ofl3_d2;
            ofl3_d4 <=  ofl3_d3;
            ofl3_d5 <=  ofl3_d4;
            ofl3_d6 <=  ofl3_d5;
            ufl2_d1 <=  ufl2;
            ufl2_d2 <=  ufl2_d1;
            ufl2_d3 <=  ufl2_d2;
            ufl2_d4 <=  ufl2_d3;
            ufl2_d5 <=  ufl2_d4;
            ufl2_d6 <=  ufl2_d5;
            ufl3_d1 <=  ufl3;
            ufl3_d2 <=  ufl3_d1;
            ufl3_d3 <=  ufl3_d2;
            ufl3_d4 <=  ufl3_d3;
            ufl3_d5 <=  ufl3_d4;
         end if;
      end process;
   Xexn <= X(wE+wFIn+2 downto wE+wFIn+1);
   XSign <= X(wE+wFIn);
   XexpField <= X(wE+wFIn-1 downto wFIn);
   Xfrac <= unsigned(X(wFIn-1 downto 0));
   e0 <= conv_std_logic_vector(113, wE+2);  -- bias - (wF+g)
   shiftVal <= ("00" & XexpField) - e0; -- for a left shift
   -- underflow when input is shifted to zero (shiftval<0), in which case exp = 1
   resultWillBeOne <= shiftVal(wE+1);
   --  mantissa with implicit bit
   mXu <= "1" & Xfrac;
   -- Partial overflow detection
   maxShift <= conv_std_logic_vector(20, wE+1);  -- wE-2 + wF+g
   overflow0 <= not shiftVal_d1(wE+1) when shiftVal_d1(wE downto 0) > maxShift_d1 else '0';
   shiftValIn <= shiftVal(4 downto 0);
   mantissa_shift: LeftShifter11_by_max_20_Freq500_uid4
      port map ( clk  => clk,
                 S => shiftValIn,
                 X => std_logic_vector(mXu),
                 R => fixX0);
   ufixX <=  unsigned(fixX0(30 downto 10)) when resultWillBeOne_d1='0' else "000000000000000000000";
   exp_helper: Exp_8_10_Freq500_uid6
      port map ( clk  => clk,
                 XSign => XSign,
                 ufixX_i => std_logic_vector(ufixX),
                 K => K,
                 expY => expY);
   needNoNorm <= expY(14);
   -- Rounding: all this should consume one row of LUTs
   preRoundBiasSig <= conv_std_logic_vector(127, wE+2)  & expY(13 downto 4) when needNoNorm = '1'
      else conv_std_logic_vector(126, wE+2)  & expY(12 downto 3) ;
   roundBit <= expY(3)  when needNoNorm = '1'    else expY(2) ;
   roundNormAddend <= K_d2(8) & K_d2 & (9 downto 1 => '0') & roundBit;
   roundedExpSigOperandAdder: IntAdder_20_Freq500_uid52
      port map ( clk  => clk,
                 Cin => '0',
                 X => preRoundBiasSig,
                 Y => roundNormAddend,
                 R => roundedExpSigRes);
   roundedExpSig <= roundedExpSigRes when Xexn_d6="01" else  "000" & (wE-2 downto 0 => '1') & (wF-1 downto 0 => '0');
   ofl1 <= not XSign_d1 and overflow0 and (not Xexn_d1(1) and Xexn_d1(0)); -- input positive, normal,  very large
   ofl2 <= not XSign_d6 and (roundedExpSig(wE+wF) and not roundedExpSig(wE+wF+1)) and (not Xexn_d6(1) and Xexn_d6(0)); -- input positive, normal, overflowed
   ofl3 <= not XSign and Xexn(1) and not Xexn(0);  -- input was -infty
   ofl <= ofl1_d5 or ofl2 or ofl3_d6;
   ufl1 <= (roundedExpSig(wE+wF) and roundedExpSig(wE+wF+1))  and (not Xexn_d6(1) and Xexn_d6(0)); -- input normal
   ufl2 <= XSign and Xexn(1) and not Xexn(0);  -- input was -infty
   ufl3 <= XSign_d1 and overflow0  and (not Xexn_d1(1) and Xexn_d1(0)); -- input negative, normal,  very large
   ufl <= ufl1 or ufl2_d6 or ufl3_d5;
   Rexn <= "11" when Xexn_d6 = "11"
      else "10" when ofl='1'
      else "00" when ufl='1'
      else "01";
   R <= Rexn & '0' & roundedExpSig(17 downto 0);
end architecture;

--------------------------------------------------------------------------------
--                     TestBench_top_module_Freq500_uid54
-- VHDL generated for DummyFPGA @ 500MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Cristian Klein, Nicolas Brunie (2007-2010)
--------------------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity TestBench_top_module_Freq500_uid54 is
end entity;

architecture behavorial of TestBench_top_module_Freq500_uid54 is
   component top_module is
      port ( clk : in std_logic;
             X : in  std_logic_vector(8+10+2 downto 0);
             R : out  std_logic_vector(8+10+2 downto 0)   );
   end component;
signal X :  std_logic_vector(20 downto 0);
   -- timing of X: (c0, 0.000000ns)
signal R :  std_logic_vector(20 downto 0);
   -- timing of R: (c6, 0.000000ns)
signal clk :  std_logic;
   -- timing of clk: (c0, 0.000000ns)
signal rst :  std_logic;
   -- timing of rst: (c0, 0.000000ns)

 -- converts std_logic into a character
   function chr(sl: std_logic) return character is
      variable c: character;
   begin
      case sl is
         when 'U' => c:= 'U';
         when 'X' => c:= 'X';
         when '0' => c:= '0';
         when '1' => c:= '1';
         when 'Z' => c:= 'Z';
         when 'W' => c:= 'W';
         when 'L' => c:= 'L';
         when 'H' => c:= 'H';
         when '-' => c:= '-';
      end case;
      return c;
   end chr;

   -- converts bit to std_logic (1 to 1)
   function to_stdlogic(b : bit) return std_logic is
       variable sl : std_logic;
   begin
      case b is 
         when '0' => sl := '0';
         when '1' => sl := '1';
      end case;
      return sl;
   end to_stdlogic;

   -- converts std_logic into a string (1 to 1)
   function str(sl: std_logic) return string is
    variable s: string(1 to 1);
    begin
      s(1) := chr(sl);
      return s;
   end str;

   -- converts std_logic_vector into a string (binary base)
   -- (this also takes care of the fact that the range of
   --  a string is natural while a std_logic_vector may
   --  have an integer range)
   function str(slv: std_logic_vector) return string is
      variable result : string (1 to slv'length);
      variable r : integer;
   begin
      r := 1;
      for i in slv'range loop
         result(r) := chr(slv(i));
         r := r + 1;
      end loop;
      return result;
   end str;

   -- FP compare function (found vs. real)
   function fp_equal(a : std_logic_vector; b : std_logic_vector) return boolean is
   begin
      if b(b'high downto b'high-1) = "01" then
         return a = b;
      elsif b(b'high downto b'high-1) = "11" then
         return (a(a'high downto a'high-1)=b(b'high downto b'high-1));
      else
         return a(a'high downto a'high-2) = b(b'high downto b'high-2);
      end if;
   end;

   function fp_inf_or_equal(a : std_logic_vector; b : std_logic_vector) return boolean is
   begin
      if (b(b'high downto b'high-1) = "11") or (a(a'high downto a'high-1) = "11")  then
         return false; -- NaN always compare false
      else return true; -- TODO
      end if;
   end;

   -- FP subtypes for casting
   subtype fp21 is std_logic_vector(20 downto 0);
   function testLine(testCounter:integer; expectedOutputS: string(1 to 10000); expectedOutputSize: integer; R:  std_logic_vector(8+10+2 downto 0)) return boolean is
      variable expectedOutput: line;
      variable possibilityNumber : integer;
      variable testSuccess: boolean;
      variable errorMessage: string(1 to 10000);
      variable testSuccess_R: boolean;
      variable expected_R: bit_vector (20 downto 0); -- for list of values
      variable inf_R: bit_vector (20 downto 0); -- for intervals
      variable sup_R: bit_vector (20 downto 0); -- for intervals
   begin
      write(expectedOutput, expectedOutputS);
      read(expectedOutput, possibilityNumber); -- for R
      if possibilityNumber = 0 then
         -- TODO define what it means to have 0 possible output. Currently it means a test fails...
      end if;
      if possibilityNumber > 0 then -- a list of values
      testSuccess_R := false;
         for i in 1 to possibilityNumber loop
            read(expectedOutput, expected_R);
            if fp_equal(R, to_stdlogicvector(expected_R)) then
               testSuccess_R := true;
            end if;
            end loop;
      end if;
      if possibilityNumber < 0  then -- an interval
         read(expectedOutput, inf_R);
         read(expectedOutput, sup_R);
         if possibilityNumber =-1  then -- an unsigned interval
            testSuccess_R := (R >= to_stdlogicvector(inf_R)) and (R <= to_stdlogicvector(sup_R));
         elsif possibilityNumber =-2  then -- a signed interval
            testSuccess_R := (signed(R) >= signed(to_stdlogicvector(inf_R))) and (signed(R) <= signed(to_stdlogicvector(sup_R)));
         elsif possibilityNumber =-4  then -- a floating-point interval
            testSuccess_R := fp_inf_or_equal(to_stdlogicvector(inf_R), R) and fp_inf_or_equal(R, to_stdlogicvector(sup_R));
         end if;
      end if;
      if testSuccess_R = false then
         report("Test #" & integer'image(testCounter) & ", incorrect output for R: " & lf & " expected values: " & expectedOutputS(1 to expectedOutputSize) & lf  & "          result:    " & str(R) ) severity error;
      end if;
      
      testSuccess := true and testSuccess_R;
      return testSuccess;
   end testLine;

begin
   -- Ticking clock signal
   process
   begin
      clk <= '0';
      wait for 5 ns;
      clk <= '1';
      wait for 5 ns;
   end process;

   test: top_module
      port map ( clk  => clk,
                 X => X,
                 R => R);
   -- Process that sets the inputs  (read from a file) 
   process
      variable input, expectedOutput : line; 
      variable tmpChar : character;
      file inputsFile : text is "test.input"; 
      variable V_X : bit_vector(20 downto 0);
      variable V_R : bit_vector(20 downto 0);
   begin
      -- Send reset
      rst <= '1';
      wait for 10 ns;
      rst <= '0';
      readline(inputsFile, input); -- skip the first line of advertising
      while not endfile(inputsFile) loop
         readline(inputsFile, input); -- skip the comment line
         readline(inputsFile, input);
         readline(inputsFile, expectedOutput); -- comment line, unused in this process
         readline(inputsFile, expectedOutput); -- unused in this process
         read(input ,V_X);
         read(input,tmpChar);
         X <= to_stdlogicvector(V_X);
         wait for 10 ns;
      end loop;
         wait for 160 ns; -- wait for pipeline to flush (and some more)
   end process;

    -- Process that verifies the corresponding output
   process
      file inputsFile : text is "test.input"; 
      variable input, expectedOutput : line; 
      variable testCounter : integer := 1;
      variable errorCounter : integer := 0;
      variable expectedOutputString : string(1 to 10000);
      variable testSuccess: boolean;
   begin
      wait for 12 ns; -- wait for reset 
      wait for 60 ns; -- wait for pipeline to flush
      readline(inputsFile, input); -- skip the first line of advertising
      while not endfile(inputsFile) loop
         readline(inputsFile, input); -- input comment, unused
         readline(inputsFile, input); -- input line, unused
         readline(inputsFile, expectedOutput); -- comment line, unused in this process
         readline(inputsFile, expectedOutput);
         expectedOutputString := expectedOutput.all & (expectedOutput'Length+1 to 10000 => ' ');
         testSuccess := testLine(testCounter, expectedOutputString, expectedOutput'Length, R);
         if not testSuccess then 
               errorCounter := errorCounter + 1; -- incrementing global error counter
         end if;
            testCounter := testCounter + 1; -- incrementing global error counter
         wait for 10 ns;
      end loop;
      report integer'image(errorCounter) & " error(s) encoutered." severity note;
      report "End of simulation after " & integer'image(testCounter-1) & " tests" severity note;
   end process;

end architecture;

