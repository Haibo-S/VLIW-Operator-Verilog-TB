module intadder_17_freq500_uid30
  (input  clk,
   input  [16:0] x,
   input  [16:0] y,
   input  cin,
   output [16:0] r);
  wire [16:0] rtmp;
  wire [16:0] x_d1;
  wire [16:0] y_d1;
  wire cin_d1;
  wire cin_d2;
  wire cin_d3;
  wire [16:0] n2259;
  wire [16:0] n2260;
  wire [16:0] n2261;
  reg [16:0] n2262;
  reg [16:0] n2263;
  reg n2264;
  reg n2265;
  reg n2266;
  assign r = rtmp; //(module output)
  /* fpexpbf16.vhdl:1132:8  */
  assign rtmp = n2261; // (signal)
  /* fpexpbf16.vhdl:1134:8  */
  assign x_d1 = n2262; // (signal)
  /* fpexpbf16.vhdl:1136:8  */
  assign y_d1 = n2263; // (signal)
  /* fpexpbf16.vhdl:1138:8  */
  assign cin_d1 = n2264; // (signal)
  /* fpexpbf16.vhdl:1138:16  */
  assign cin_d2 = n2265; // (signal)
  /* fpexpbf16.vhdl:1138:24  */
  assign cin_d3 = n2266; // (signal)
  /* fpexpbf16.vhdl:1151:17  */
  assign n2259 = x_d1 + y_d1;
  /* fpexpbf16.vhdl:1151:24  */
  assign n2260 = {16'b0, cin_d3};  //  uext
  /* fpexpbf16.vhdl:1151:24  */
  assign n2261 = n2259 + n2260;
  /* fpexpbf16.vhdl:1143:10  */
  always @(posedge clk)
    n2262 <= x;
  /* fpexpbf16.vhdl:1143:10  */
  always @(posedge clk)
    n2263 <= y;
  /* fpexpbf16.vhdl:1143:10  */
  always @(posedge clk)
    n2264 <= cin;
  /* fpexpbf16.vhdl:1143:10  */
  always @(posedge clk)
    n2265 <= cin_d1;
  /* fpexpbf16.vhdl:1143:10  */
  always @(posedge clk)
    n2266 <= cin_d2;
endmodule

module fixrealkcm_freq500_uid20_t1_freq500_uid26
  (input  [2:0] x,
   output [11:0] y);
  wire [11:0] y0;
  wire [11:0] y1;
  wire n2224;
  wire n2227;
  wire n2230;
  wire n2233;
  wire n2236;
  wire n2239;
  wire n2242;
  wire n2245;
  wire [7:0] n2247;
  reg [11:0] n2248;
  assign y = y1; //(module output)
  /* fpexpbf16.vhdl:246:8  */
  assign y0 = n2248; // (signal)
  /* fpexpbf16.vhdl:248:8  */
  assign y1 = y0; // (signal)
  /* fpexpbf16.vhdl:252:22  */
  assign n2224 = x == 3'b000;
  /* fpexpbf16.vhdl:253:22  */
  assign n2227 = x == 3'b001;
  /* fpexpbf16.vhdl:254:22  */
  assign n2230 = x == 3'b010;
  /* fpexpbf16.vhdl:255:22  */
  assign n2233 = x == 3'b011;
  /* fpexpbf16.vhdl:256:22  */
  assign n2236 = x == 3'b100;
  /* fpexpbf16.vhdl:257:22  */
  assign n2239 = x == 3'b101;
  /* fpexpbf16.vhdl:258:22  */
  assign n2242 = x == 3'b110;
  /* fpexpbf16.vhdl:259:22  */
  assign n2245 = x == 3'b111;
  assign n2247 = {n2245, n2242, n2239, n2236, n2233, n2230, n2227, n2224};
  /* fpexpbf16.vhdl:251:4  */
  always @*
    case (n2247)
      8'b10000000: n2248 = 12'b100110110100;
      8'b01000000: n2248 = 12'b100001010001;
      8'b00100000: n2248 = 12'b011011101110;
      8'b00010000: n2248 = 12'b010110001100;
      8'b00001000: n2248 = 12'b010000101001;
      8'b00000100: n2248 = 12'b001011000110;
      8'b00000010: n2248 = 12'b000101100011;
      8'b00000001: n2248 = 12'b000000000000;
      default: n2248 = 12'bX;
    endcase
endmodule

module fixrealkcm_freq500_uid20_t0_freq500_uid23
  (input  [4:0] x,
   output [16:0] y);
  wire [16:0] y0;
  wire [16:0] y1;
  wire n2124;
  wire n2127;
  wire n2130;
  wire n2133;
  wire n2136;
  wire n2139;
  wire n2142;
  wire n2145;
  wire n2148;
  wire n2151;
  wire n2154;
  wire n2157;
  wire n2160;
  wire n2163;
  wire n2166;
  wire n2169;
  wire n2172;
  wire n2175;
  wire n2178;
  wire n2181;
  wire n2184;
  wire n2187;
  wire n2190;
  wire n2193;
  wire n2196;
  wire n2199;
  wire n2202;
  wire n2205;
  wire n2208;
  wire n2211;
  wire n2214;
  wire n2217;
  wire [31:0] n2219;
  reg [16:0] n2220;
  assign y = y1; //(module output)
  /* fpexpbf16.vhdl:174:8  */
  assign y0 = n2220; // (signal)
  /* fpexpbf16.vhdl:176:8  */
  assign y1 = y0; // (signal)
  /* fpexpbf16.vhdl:180:27  */
  assign n2124 = x == 5'b00000;
  /* fpexpbf16.vhdl:181:27  */
  assign n2127 = x == 5'b00001;
  /* fpexpbf16.vhdl:182:27  */
  assign n2130 = x == 5'b00010;
  /* fpexpbf16.vhdl:183:27  */
  assign n2133 = x == 5'b00011;
  /* fpexpbf16.vhdl:184:27  */
  assign n2136 = x == 5'b00100;
  /* fpexpbf16.vhdl:185:27  */
  assign n2139 = x == 5'b00101;
  /* fpexpbf16.vhdl:186:27  */
  assign n2142 = x == 5'b00110;
  /* fpexpbf16.vhdl:187:27  */
  assign n2145 = x == 5'b00111;
  /* fpexpbf16.vhdl:188:27  */
  assign n2148 = x == 5'b01000;
  /* fpexpbf16.vhdl:189:27  */
  assign n2151 = x == 5'b01001;
  /* fpexpbf16.vhdl:190:27  */
  assign n2154 = x == 5'b01010;
  /* fpexpbf16.vhdl:191:27  */
  assign n2157 = x == 5'b01011;
  /* fpexpbf16.vhdl:192:27  */
  assign n2160 = x == 5'b01100;
  /* fpexpbf16.vhdl:193:27  */
  assign n2163 = x == 5'b01101;
  /* fpexpbf16.vhdl:194:27  */
  assign n2166 = x == 5'b01110;
  /* fpexpbf16.vhdl:195:27  */
  assign n2169 = x == 5'b01111;
  /* fpexpbf16.vhdl:196:27  */
  assign n2172 = x == 5'b10000;
  /* fpexpbf16.vhdl:197:27  */
  assign n2175 = x == 5'b10001;
  /* fpexpbf16.vhdl:198:27  */
  assign n2178 = x == 5'b10010;
  /* fpexpbf16.vhdl:199:27  */
  assign n2181 = x == 5'b10011;
  /* fpexpbf16.vhdl:200:27  */
  assign n2184 = x == 5'b10100;
  /* fpexpbf16.vhdl:201:27  */
  assign n2187 = x == 5'b10101;
  /* fpexpbf16.vhdl:202:27  */
  assign n2190 = x == 5'b10110;
  /* fpexpbf16.vhdl:203:27  */
  assign n2193 = x == 5'b10111;
  /* fpexpbf16.vhdl:204:27  */
  assign n2196 = x == 5'b11000;
  /* fpexpbf16.vhdl:205:27  */
  assign n2199 = x == 5'b11001;
  /* fpexpbf16.vhdl:206:27  */
  assign n2202 = x == 5'b11010;
  /* fpexpbf16.vhdl:207:27  */
  assign n2205 = x == 5'b11011;
  /* fpexpbf16.vhdl:208:27  */
  assign n2208 = x == 5'b11100;
  /* fpexpbf16.vhdl:209:27  */
  assign n2211 = x == 5'b11101;
  /* fpexpbf16.vhdl:210:27  */
  assign n2214 = x == 5'b11110;
  /* fpexpbf16.vhdl:211:27  */
  assign n2217 = x == 5'b11111;
  assign n2219 = {n2217, n2214, n2211, n2208, n2205, n2202, n2199, n2196, n2193, n2190, n2187, n2184, n2181, n2178, n2175, n2172, n2169, n2166, n2163, n2160, n2157, n2154, n2151, n2148, n2145, n2142, n2139, n2136, n2133, n2130, n2127, n2124};
  /* fpexpbf16.vhdl:179:4  */
  always @*
    case (n2219)
      32'b10000000000000000000000000000000: n2220 = 17'b10101011111001101;
      32'b01000000000000000000000000000000: n2220 = 17'b10100110010110110;
      32'b00100000000000000000000000000000: n2220 = 17'b10100000110011111;
      32'b00010000000000000000000000000000: n2220 = 17'b10011011010001000;
      32'b00001000000000000000000000000000: n2220 = 17'b10010101101110001;
      32'b00000100000000000000000000000000: n2220 = 17'b10010000001011001;
      32'b00000010000000000000000000000000: n2220 = 17'b10001010101000010;
      32'b00000001000000000000000000000000: n2220 = 17'b10000101000101011;
      32'b00000000100000000000000000000000: n2220 = 17'b01111111100010100;
      32'b00000000010000000000000000000000: n2220 = 17'b01111001111111101;
      32'b00000000001000000000000000000000: n2220 = 17'b01110100011100110;
      32'b00000000000100000000000000000000: n2220 = 17'b01101110111001111;
      32'b00000000000010000000000000000000: n2220 = 17'b01101001010110111;
      32'b00000000000001000000000000000000: n2220 = 17'b01100011110100000;
      32'b00000000000000100000000000000000: n2220 = 17'b01011110010001001;
      32'b00000000000000010000000000000000: n2220 = 17'b01011000101110010;
      32'b00000000000000001000000000000000: n2220 = 17'b01010011001011011;
      32'b00000000000000000100000000000000: n2220 = 17'b01001101101000100;
      32'b00000000000000000010000000000000: n2220 = 17'b01001000000101101;
      32'b00000000000000000001000000000000: n2220 = 17'b01000010100010110;
      32'b00000000000000000000100000000000: n2220 = 17'b00111100111111110;
      32'b00000000000000000000010000000000: n2220 = 17'b00110111011100111;
      32'b00000000000000000000001000000000: n2220 = 17'b00110001111010000;
      32'b00000000000000000000000100000000: n2220 = 17'b00101100010111001;
      32'b00000000000000000000000010000000: n2220 = 17'b00100110110100010;
      32'b00000000000000000000000001000000: n2220 = 17'b00100001010001011;
      32'b00000000000000000000000000100000: n2220 = 17'b00011011101110100;
      32'b00000000000000000000000000010000: n2220 = 17'b00010110001011101;
      32'b00000000000000000000000000001000: n2220 = 17'b00010000101000101;
      32'b00000000000000000000000000000100: n2220 = 17'b00001011000101110;
      32'b00000000000000000000000000000010: n2220 = 17'b00000101100010111;
      32'b00000000000000000000000000000001: n2220 = 17'b00000000000000000;
      default: n2220 = 17'bX;
    endcase
endmodule

module intadder_12_freq500_uid18
  (input  clk,
   input  [11:0] x,
   input  [11:0] y,
   input  cin,
   output [11:0] r);
  wire cin_1;
  wire cin_1_d1;
  wire cin_1_d2;
  wire [12:0] x_1;
  wire [12:0] x_1_d1;
  wire [12:0] y_1;
  wire [12:0] y_1_d1;
  wire [12:0] s_1;
  wire [11:0] r_1;
  wire [12:0] n2110;
  wire [12:0] n2112;
  wire [12:0] n2113;
  wire [12:0] n2114;
  wire [12:0] n2115;
  wire [11:0] n2116;
  reg n2117;
  reg n2118;
  reg [12:0] n2119;
  reg [12:0] n2120;
  assign r = r_1; //(module output)
  /* fpexpbf16.vhdl:911:15  */
  assign cin_1_d1 = n2117; // (signal)
  /* fpexpbf16.vhdl:911:25  */
  assign cin_1_d2 = n2118; // (signal)
  /* fpexpbf16.vhdl:913:8  */
  assign x_1 = n2110; // (signal)
  /* fpexpbf16.vhdl:913:13  */
  assign x_1_d1 = n2119; // (signal)
  /* fpexpbf16.vhdl:915:8  */
  assign y_1 = n2112; // (signal)
  /* fpexpbf16.vhdl:915:13  */
  assign y_1_d1 = n2120; // (signal)
  /* fpexpbf16.vhdl:917:8  */
  assign s_1 = n2115; // (signal)
  /* fpexpbf16.vhdl:919:8  */
  assign r_1 = n2116; // (signal)
  /* fpexpbf16.vhdl:932:15  */
  assign n2110 = {1'b0, x};
  /* fpexpbf16.vhdl:933:15  */
  assign n2112 = {1'b0, y};
  /* fpexpbf16.vhdl:934:18  */
  assign n2113 = x_1_d1 + y_1_d1;
  /* fpexpbf16.vhdl:934:27  */
  assign n2114 = {12'b0, cin_1_d2};  //  uext
  /* fpexpbf16.vhdl:934:27  */
  assign n2115 = n2113 + n2114;
  /* fpexpbf16.vhdl:935:14  */
  assign n2116 = s_1[11:0]; // extract
  /* fpexpbf16.vhdl:924:10  */
  always @(posedge clk)
    n2117 <= cin_1;
  /* fpexpbf16.vhdl:924:10  */
  always @(posedge clk)
    n2118 <= cin_1_d1;
  /* fpexpbf16.vhdl:924:10  */
  always @(posedge clk)
    n2119 <= x_1;
  /* fpexpbf16.vhdl:924:10  */
  always @(posedge clk)
    n2120 <= y_1;
endmodule

module fixrealkcm_freq500_uid8_t1_freq500_uid14
  (input  [4:0] x,
   output [6:0] y);
  wire [6:0] y0;
  wire [6:0] y1;
  wire n2003;
  wire n2006;
  wire n2009;
  wire n2012;
  wire n2015;
  wire n2018;
  wire n2021;
  wire n2024;
  wire n2027;
  wire n2030;
  wire n2033;
  wire n2036;
  wire n2039;
  wire n2042;
  wire n2045;
  wire n2048;
  wire n2051;
  wire n2054;
  wire n2057;
  wire n2060;
  wire n2063;
  wire n2066;
  wire n2069;
  wire n2072;
  wire n2075;
  wire n2078;
  wire n2081;
  wire n2084;
  wire n2087;
  wire n2090;
  wire n2093;
  wire n2096;
  wire [31:0] n2098;
  reg [6:0] n2099;
  assign y = y1; //(module output)
  /* fpexpbf16.vhdl:102:8  */
  assign y0 = n2099; // (signal)
  /* fpexpbf16.vhdl:104:8  */
  assign y1 = y0; // (signal)
  /* fpexpbf16.vhdl:108:17  */
  assign n2003 = x == 5'b00000;
  /* fpexpbf16.vhdl:109:17  */
  assign n2006 = x == 5'b00001;
  /* fpexpbf16.vhdl:110:17  */
  assign n2009 = x == 5'b00010;
  /* fpexpbf16.vhdl:111:17  */
  assign n2012 = x == 5'b00011;
  /* fpexpbf16.vhdl:112:17  */
  assign n2015 = x == 5'b00100;
  /* fpexpbf16.vhdl:113:17  */
  assign n2018 = x == 5'b00101;
  /* fpexpbf16.vhdl:114:17  */
  assign n2021 = x == 5'b00110;
  /* fpexpbf16.vhdl:115:17  */
  assign n2024 = x == 5'b00111;
  /* fpexpbf16.vhdl:116:17  */
  assign n2027 = x == 5'b01000;
  /* fpexpbf16.vhdl:117:17  */
  assign n2030 = x == 5'b01001;
  /* fpexpbf16.vhdl:118:17  */
  assign n2033 = x == 5'b01010;
  /* fpexpbf16.vhdl:119:17  */
  assign n2036 = x == 5'b01011;
  /* fpexpbf16.vhdl:120:17  */
  assign n2039 = x == 5'b01100;
  /* fpexpbf16.vhdl:121:17  */
  assign n2042 = x == 5'b01101;
  /* fpexpbf16.vhdl:122:17  */
  assign n2045 = x == 5'b01110;
  /* fpexpbf16.vhdl:123:17  */
  assign n2048 = x == 5'b01111;
  /* fpexpbf16.vhdl:124:17  */
  assign n2051 = x == 5'b10000;
  /* fpexpbf16.vhdl:125:17  */
  assign n2054 = x == 5'b10001;
  /* fpexpbf16.vhdl:126:17  */
  assign n2057 = x == 5'b10010;
  /* fpexpbf16.vhdl:127:17  */
  assign n2060 = x == 5'b10011;
  /* fpexpbf16.vhdl:128:17  */
  assign n2063 = x == 5'b10100;
  /* fpexpbf16.vhdl:129:17  */
  assign n2066 = x == 5'b10101;
  /* fpexpbf16.vhdl:130:17  */
  assign n2069 = x == 5'b10110;
  /* fpexpbf16.vhdl:131:17  */
  assign n2072 = x == 5'b10111;
  /* fpexpbf16.vhdl:132:17  */
  assign n2075 = x == 5'b11000;
  /* fpexpbf16.vhdl:133:17  */
  assign n2078 = x == 5'b11001;
  /* fpexpbf16.vhdl:134:17  */
  assign n2081 = x == 5'b11010;
  /* fpexpbf16.vhdl:135:17  */
  assign n2084 = x == 5'b11011;
  /* fpexpbf16.vhdl:136:17  */
  assign n2087 = x == 5'b11100;
  /* fpexpbf16.vhdl:137:17  */
  assign n2090 = x == 5'b11101;
  /* fpexpbf16.vhdl:138:17  */
  assign n2093 = x == 5'b11110;
  /* fpexpbf16.vhdl:139:17  */
  assign n2096 = x == 5'b11111;
  assign n2098 = {n2096, n2093, n2090, n2087, n2084, n2081, n2078, n2075, n2072, n2069, n2066, n2063, n2060, n2057, n2054, n2051, n2048, n2045, n2042, n2039, n2036, n2033, n2030, n2027, n2024, n2021, n2018, n2015, n2012, n2009, n2006, n2003};
  /* fpexpbf16.vhdl:107:4  */
  always @*
    case (n2098)
      32'b10000000000000000000000000000000: n2099 = 7'b1011001;
      32'b01000000000000000000000000000000: n2099 = 7'b1010111;
      32'b00100000000000000000000000000000: n2099 = 7'b1010100;
      32'b00010000000000000000000000000000: n2099 = 7'b1010001;
      32'b00001000000000000000000000000000: n2099 = 7'b1001110;
      32'b00000100000000000000000000000000: n2099 = 7'b1001011;
      32'b00000010000000000000000000000000: n2099 = 7'b1001000;
      32'b00000001000000000000000000000000: n2099 = 7'b1000101;
      32'b00000000100000000000000000000000: n2099 = 7'b1000010;
      32'b00000000010000000000000000000000: n2099 = 7'b0111111;
      32'b00000000001000000000000000000000: n2099 = 7'b0111101;
      32'b00000000000100000000000000000000: n2099 = 7'b0111010;
      32'b00000000000010000000000000000000: n2099 = 7'b0110111;
      32'b00000000000001000000000000000000: n2099 = 7'b0110100;
      32'b00000000000000100000000000000000: n2099 = 7'b0110001;
      32'b00000000000000010000000000000000: n2099 = 7'b0101110;
      32'b00000000000000001000000000000000: n2099 = 7'b0101011;
      32'b00000000000000000100000000000000: n2099 = 7'b0101000;
      32'b00000000000000000010000000000000: n2099 = 7'b0100110;
      32'b00000000000000000001000000000000: n2099 = 7'b0100011;
      32'b00000000000000000000100000000000: n2099 = 7'b0100000;
      32'b00000000000000000000010000000000: n2099 = 7'b0011101;
      32'b00000000000000000000001000000000: n2099 = 7'b0011010;
      32'b00000000000000000000000100000000: n2099 = 7'b0010111;
      32'b00000000000000000000000010000000: n2099 = 7'b0010100;
      32'b00000000000000000000000001000000: n2099 = 7'b0010001;
      32'b00000000000000000000000000100000: n2099 = 7'b0001110;
      32'b00000000000000000000000000010000: n2099 = 7'b0001100;
      32'b00000000000000000000000000001000: n2099 = 7'b0001001;
      32'b00000000000000000000000000000100: n2099 = 7'b0000110;
      32'b00000000000000000000000000000010: n2099 = 7'b0000011;
      32'b00000000000000000000000000000001: n2099 = 7'b0000000;
      default: n2099 = 7'bX;
    endcase
endmodule

module fixrealkcm_freq500_uid8_t0_freq500_uid11
  (input  [4:0] x,
   output [11:0] y);
  wire [11:0] y0;
  wire [11:0] y1;
  wire n1903;
  wire n1906;
  wire n1909;
  wire n1912;
  wire n1915;
  wire n1918;
  wire n1921;
  wire n1924;
  wire n1927;
  wire n1930;
  wire n1933;
  wire n1936;
  wire n1939;
  wire n1942;
  wire n1945;
  wire n1948;
  wire n1951;
  wire n1954;
  wire n1957;
  wire n1960;
  wire n1963;
  wire n1966;
  wire n1969;
  wire n1972;
  wire n1975;
  wire n1978;
  wire n1981;
  wire n1984;
  wire n1987;
  wire n1990;
  wire n1993;
  wire n1996;
  wire [31:0] n1998;
  reg [11:0] n1999;
  assign y = y1; //(module output)
  /* fpexpbf16.vhdl:30:8  */
  assign y0 = n1999; // (signal)
  /* fpexpbf16.vhdl:32:8  */
  assign y1 = y0; // (signal)
  /* fpexpbf16.vhdl:36:22  */
  assign n1903 = x == 5'b00000;
  /* fpexpbf16.vhdl:37:22  */
  assign n1906 = x == 5'b00001;
  /* fpexpbf16.vhdl:38:22  */
  assign n1909 = x == 5'b00010;
  /* fpexpbf16.vhdl:39:22  */
  assign n1912 = x == 5'b00011;
  /* fpexpbf16.vhdl:40:22  */
  assign n1915 = x == 5'b00100;
  /* fpexpbf16.vhdl:41:22  */
  assign n1918 = x == 5'b00101;
  /* fpexpbf16.vhdl:42:22  */
  assign n1921 = x == 5'b00110;
  /* fpexpbf16.vhdl:43:22  */
  assign n1924 = x == 5'b00111;
  /* fpexpbf16.vhdl:44:22  */
  assign n1927 = x == 5'b01000;
  /* fpexpbf16.vhdl:45:22  */
  assign n1930 = x == 5'b01001;
  /* fpexpbf16.vhdl:46:22  */
  assign n1933 = x == 5'b01010;
  /* fpexpbf16.vhdl:47:22  */
  assign n1936 = x == 5'b01011;
  /* fpexpbf16.vhdl:48:22  */
  assign n1939 = x == 5'b01100;
  /* fpexpbf16.vhdl:49:22  */
  assign n1942 = x == 5'b01101;
  /* fpexpbf16.vhdl:50:22  */
  assign n1945 = x == 5'b01110;
  /* fpexpbf16.vhdl:51:22  */
  assign n1948 = x == 5'b01111;
  /* fpexpbf16.vhdl:52:22  */
  assign n1951 = x == 5'b10000;
  /* fpexpbf16.vhdl:53:22  */
  assign n1954 = x == 5'b10001;
  /* fpexpbf16.vhdl:54:22  */
  assign n1957 = x == 5'b10010;
  /* fpexpbf16.vhdl:55:22  */
  assign n1960 = x == 5'b10011;
  /* fpexpbf16.vhdl:56:22  */
  assign n1963 = x == 5'b10100;
  /* fpexpbf16.vhdl:57:22  */
  assign n1966 = x == 5'b10101;
  /* fpexpbf16.vhdl:58:22  */
  assign n1969 = x == 5'b10110;
  /* fpexpbf16.vhdl:59:22  */
  assign n1972 = x == 5'b10111;
  /* fpexpbf16.vhdl:60:22  */
  assign n1975 = x == 5'b11000;
  /* fpexpbf16.vhdl:61:22  */
  assign n1978 = x == 5'b11001;
  /* fpexpbf16.vhdl:62:22  */
  assign n1981 = x == 5'b11010;
  /* fpexpbf16.vhdl:63:22  */
  assign n1984 = x == 5'b11011;
  /* fpexpbf16.vhdl:64:22  */
  assign n1987 = x == 5'b11100;
  /* fpexpbf16.vhdl:65:22  */
  assign n1990 = x == 5'b11101;
  /* fpexpbf16.vhdl:66:22  */
  assign n1993 = x == 5'b11110;
  /* fpexpbf16.vhdl:67:22  */
  assign n1996 = x == 5'b11111;
  assign n1998 = {n1996, n1993, n1990, n1987, n1984, n1981, n1978, n1975, n1972, n1969, n1966, n1963, n1960, n1957, n1954, n1951, n1948, n1945, n1942, n1939, n1936, n1933, n1930, n1927, n1924, n1921, n1918, n1915, n1912, n1909, n1906, n1903};
  /* fpexpbf16.vhdl:35:4  */
  always @*
    case (n1998)
      32'b10000000000000000000000000000000: n1999 = 12'b101100110110;
      32'b01000000000000000000000000000000: n1999 = 12'b101011011010;
      32'b00100000000000000000000000000000: n1999 = 12'b101001111110;
      32'b00010000000000000000000000000000: n1999 = 12'b101000100001;
      32'b00001000000000000000000000000000: n1999 = 12'b100111000101;
      32'b00000100000000000000000000000000: n1999 = 12'b100101101001;
      32'b00000010000000000000000000000000: n1999 = 12'b100100001100;
      32'b00000001000000000000000000000000: n1999 = 12'b100010110000;
      32'b00000000100000000000000000000000: n1999 = 12'b100001010100;
      32'b00000000010000000000000000000000: n1999 = 12'b011111110111;
      32'b00000000001000000000000000000000: n1999 = 12'b011110011011;
      32'b00000000000100000000000000000000: n1999 = 12'b011100111111;
      32'b00000000000010000000000000000000: n1999 = 12'b011011100010;
      32'b00000000000001000000000000000000: n1999 = 12'b011010000110;
      32'b00000000000000100000000000000000: n1999 = 12'b011000101010;
      32'b00000000000000010000000000000000: n1999 = 12'b010111001101;
      32'b00000000000000001000000000000000: n1999 = 12'b010101110001;
      32'b00000000000000000100000000000000: n1999 = 12'b010100010101;
      32'b00000000000000000010000000000000: n1999 = 12'b010010111000;
      32'b00000000000000000001000000000000: n1999 = 12'b010001011100;
      32'b00000000000000000000100000000000: n1999 = 12'b010000000000;
      32'b00000000000000000000010000000000: n1999 = 12'b001110100011;
      32'b00000000000000000000001000000000: n1999 = 12'b001101000111;
      32'b00000000000000000000000100000000: n1999 = 12'b001011101011;
      32'b00000000000000000000000010000000: n1999 = 12'b001010001110;
      32'b00000000000000000000000001000000: n1999 = 12'b001000110010;
      32'b00000000000000000000000000100000: n1999 = 12'b000111010110;
      32'b00000000000000000000000000010000: n1999 = 12'b000101111001;
      32'b00000000000000000000000000001000: n1999 = 12'b000100011101;
      32'b00000000000000000000000000000100: n1999 = 12'b000011000001;
      32'b00000000000000000000000000000010: n1999 = 12'b000001100100;
      32'b00000000000000000000000000000001: n1999 = 12'b000000001000;
      default: n1999 = 12'bX;
    endcase
endmodule

module fixfunctionbytable_freq500_uid35
  (input  [8:0] x,
   output [11:0] y);
  wire [11:0] y0;
  wire [11:0] y1;
  wire n363;
  wire n366;
  wire n369;
  wire n372;
  wire n375;
  wire n378;
  wire n381;
  wire n384;
  wire n387;
  wire n390;
  wire n393;
  wire n396;
  wire n399;
  wire n402;
  wire n405;
  wire n408;
  wire n411;
  wire n414;
  wire n417;
  wire n420;
  wire n423;
  wire n426;
  wire n429;
  wire n432;
  wire n435;
  wire n438;
  wire n441;
  wire n444;
  wire n447;
  wire n450;
  wire n453;
  wire n456;
  wire n459;
  wire n462;
  wire n465;
  wire n468;
  wire n471;
  wire n474;
  wire n477;
  wire n480;
  wire n483;
  wire n486;
  wire n489;
  wire n492;
  wire n495;
  wire n498;
  wire n501;
  wire n504;
  wire n507;
  wire n510;
  wire n513;
  wire n516;
  wire n519;
  wire n522;
  wire n525;
  wire n528;
  wire n531;
  wire n534;
  wire n537;
  wire n540;
  wire n543;
  wire n546;
  wire n549;
  wire n552;
  wire n555;
  wire n558;
  wire n561;
  wire n564;
  wire n567;
  wire n570;
  wire n573;
  wire n576;
  wire n579;
  wire n582;
  wire n585;
  wire n588;
  wire n591;
  wire n594;
  wire n597;
  wire n600;
  wire n603;
  wire n606;
  wire n609;
  wire n612;
  wire n615;
  wire n618;
  wire n621;
  wire n624;
  wire n627;
  wire n630;
  wire n633;
  wire n636;
  wire n639;
  wire n642;
  wire n645;
  wire n648;
  wire n651;
  wire n654;
  wire n657;
  wire n660;
  wire n663;
  wire n666;
  wire n669;
  wire n672;
  wire n675;
  wire n678;
  wire n681;
  wire n684;
  wire n687;
  wire n690;
  wire n693;
  wire n696;
  wire n699;
  wire n702;
  wire n705;
  wire n708;
  wire n711;
  wire n714;
  wire n717;
  wire n720;
  wire n723;
  wire n726;
  wire n729;
  wire n732;
  wire n735;
  wire n738;
  wire n741;
  wire n744;
  wire n747;
  wire n750;
  wire n753;
  wire n756;
  wire n759;
  wire n762;
  wire n765;
  wire n768;
  wire n771;
  wire n774;
  wire n777;
  wire n780;
  wire n783;
  wire n786;
  wire n789;
  wire n792;
  wire n795;
  wire n798;
  wire n801;
  wire n804;
  wire n807;
  wire n810;
  wire n813;
  wire n816;
  wire n819;
  wire n822;
  wire n825;
  wire n828;
  wire n831;
  wire n834;
  wire n837;
  wire n840;
  wire n843;
  wire n846;
  wire n849;
  wire n852;
  wire n855;
  wire n858;
  wire n861;
  wire n864;
  wire n867;
  wire n870;
  wire n873;
  wire n876;
  wire n879;
  wire n882;
  wire n885;
  wire n888;
  wire n891;
  wire n894;
  wire n897;
  wire n900;
  wire n903;
  wire n906;
  wire n909;
  wire n912;
  wire n915;
  wire n918;
  wire n921;
  wire n924;
  wire n927;
  wire n930;
  wire n933;
  wire n936;
  wire n939;
  wire n942;
  wire n945;
  wire n948;
  wire n951;
  wire n954;
  wire n957;
  wire n960;
  wire n963;
  wire n966;
  wire n969;
  wire n972;
  wire n975;
  wire n978;
  wire n981;
  wire n984;
  wire n987;
  wire n990;
  wire n993;
  wire n996;
  wire n999;
  wire n1002;
  wire n1005;
  wire n1008;
  wire n1011;
  wire n1014;
  wire n1017;
  wire n1020;
  wire n1023;
  wire n1026;
  wire n1029;
  wire n1032;
  wire n1035;
  wire n1038;
  wire n1041;
  wire n1044;
  wire n1047;
  wire n1050;
  wire n1053;
  wire n1056;
  wire n1059;
  wire n1062;
  wire n1065;
  wire n1068;
  wire n1071;
  wire n1074;
  wire n1077;
  wire n1080;
  wire n1083;
  wire n1086;
  wire n1089;
  wire n1092;
  wire n1095;
  wire n1098;
  wire n1101;
  wire n1104;
  wire n1107;
  wire n1110;
  wire n1113;
  wire n1116;
  wire n1119;
  wire n1122;
  wire n1125;
  wire n1128;
  wire n1131;
  wire n1134;
  wire n1137;
  wire n1140;
  wire n1143;
  wire n1146;
  wire n1149;
  wire n1152;
  wire n1155;
  wire n1158;
  wire n1161;
  wire n1164;
  wire n1167;
  wire n1170;
  wire n1173;
  wire n1176;
  wire n1179;
  wire n1182;
  wire n1185;
  wire n1188;
  wire n1191;
  wire n1194;
  wire n1197;
  wire n1200;
  wire n1203;
  wire n1206;
  wire n1209;
  wire n1212;
  wire n1215;
  wire n1218;
  wire n1221;
  wire n1224;
  wire n1227;
  wire n1230;
  wire n1233;
  wire n1236;
  wire n1239;
  wire n1242;
  wire n1245;
  wire n1248;
  wire n1251;
  wire n1254;
  wire n1257;
  wire n1260;
  wire n1263;
  wire n1266;
  wire n1269;
  wire n1272;
  wire n1275;
  wire n1278;
  wire n1281;
  wire n1284;
  wire n1287;
  wire n1290;
  wire n1293;
  wire n1296;
  wire n1299;
  wire n1302;
  wire n1305;
  wire n1308;
  wire n1311;
  wire n1314;
  wire n1317;
  wire n1320;
  wire n1323;
  wire n1326;
  wire n1329;
  wire n1332;
  wire n1335;
  wire n1338;
  wire n1341;
  wire n1344;
  wire n1347;
  wire n1350;
  wire n1353;
  wire n1356;
  wire n1359;
  wire n1362;
  wire n1365;
  wire n1368;
  wire n1371;
  wire n1374;
  wire n1377;
  wire n1380;
  wire n1383;
  wire n1386;
  wire n1389;
  wire n1392;
  wire n1395;
  wire n1398;
  wire n1401;
  wire n1404;
  wire n1407;
  wire n1410;
  wire n1413;
  wire n1416;
  wire n1419;
  wire n1422;
  wire n1425;
  wire n1428;
  wire n1431;
  wire n1434;
  wire n1437;
  wire n1440;
  wire n1443;
  wire n1446;
  wire n1449;
  wire n1452;
  wire n1455;
  wire n1458;
  wire n1461;
  wire n1464;
  wire n1467;
  wire n1470;
  wire n1473;
  wire n1476;
  wire n1479;
  wire n1482;
  wire n1485;
  wire n1488;
  wire n1491;
  wire n1494;
  wire n1497;
  wire n1500;
  wire n1503;
  wire n1506;
  wire n1509;
  wire n1512;
  wire n1515;
  wire n1518;
  wire n1521;
  wire n1524;
  wire n1527;
  wire n1530;
  wire n1533;
  wire n1536;
  wire n1539;
  wire n1542;
  wire n1545;
  wire n1548;
  wire n1551;
  wire n1554;
  wire n1557;
  wire n1560;
  wire n1563;
  wire n1566;
  wire n1569;
  wire n1572;
  wire n1575;
  wire n1578;
  wire n1581;
  wire n1584;
  wire n1587;
  wire n1590;
  wire n1593;
  wire n1596;
  wire n1599;
  wire n1602;
  wire n1605;
  wire n1608;
  wire n1611;
  wire n1614;
  wire n1617;
  wire n1620;
  wire n1623;
  wire n1626;
  wire n1629;
  wire n1632;
  wire n1635;
  wire n1638;
  wire n1641;
  wire n1644;
  wire n1647;
  wire n1650;
  wire n1653;
  wire n1656;
  wire n1659;
  wire n1662;
  wire n1665;
  wire n1668;
  wire n1671;
  wire n1674;
  wire n1677;
  wire n1680;
  wire n1683;
  wire n1686;
  wire n1689;
  wire n1692;
  wire n1695;
  wire n1698;
  wire n1701;
  wire n1704;
  wire n1707;
  wire n1710;
  wire n1713;
  wire n1716;
  wire n1719;
  wire n1722;
  wire n1725;
  wire n1728;
  wire n1731;
  wire n1734;
  wire n1737;
  wire n1740;
  wire n1743;
  wire n1746;
  wire n1749;
  wire n1752;
  wire n1755;
  wire n1758;
  wire n1761;
  wire n1764;
  wire n1767;
  wire n1770;
  wire n1773;
  wire n1776;
  wire n1779;
  wire n1782;
  wire n1785;
  wire n1788;
  wire n1791;
  wire n1794;
  wire n1797;
  wire n1800;
  wire n1803;
  wire n1806;
  wire n1809;
  wire n1812;
  wire n1815;
  wire n1818;
  wire n1821;
  wire n1824;
  wire n1827;
  wire n1830;
  wire n1833;
  wire n1836;
  wire n1839;
  wire n1842;
  wire n1845;
  wire n1848;
  wire n1851;
  wire n1854;
  wire n1857;
  wire n1860;
  wire n1863;
  wire n1866;
  wire n1869;
  wire n1872;
  wire n1875;
  wire n1878;
  wire n1881;
  wire n1884;
  wire n1887;
  wire n1890;
  wire n1893;
  wire n1896;
  wire [511:0] n1898;
  reg [11:0] n1899;
  assign y = y1; //(module output)
  /* fpexpbf16.vhdl:296:8  */
  assign y0 = n1899; // (signal)
  /* fpexpbf16.vhdl:298:8  */
  assign y1 = y0; // (signal)
  /* fpexpbf16.vhdl:302:22  */
  assign n363 = x == 9'b000000000;
  /* fpexpbf16.vhdl:303:22  */
  assign n366 = x == 9'b000000001;
  /* fpexpbf16.vhdl:304:22  */
  assign n369 = x == 9'b000000010;
  /* fpexpbf16.vhdl:305:22  */
  assign n372 = x == 9'b000000011;
  /* fpexpbf16.vhdl:306:22  */
  assign n375 = x == 9'b000000100;
  /* fpexpbf16.vhdl:307:22  */
  assign n378 = x == 9'b000000101;
  /* fpexpbf16.vhdl:308:22  */
  assign n381 = x == 9'b000000110;
  /* fpexpbf16.vhdl:309:22  */
  assign n384 = x == 9'b000000111;
  /* fpexpbf16.vhdl:310:22  */
  assign n387 = x == 9'b000001000;
  /* fpexpbf16.vhdl:311:22  */
  assign n390 = x == 9'b000001001;
  /* fpexpbf16.vhdl:312:22  */
  assign n393 = x == 9'b000001010;
  /* fpexpbf16.vhdl:313:22  */
  assign n396 = x == 9'b000001011;
  /* fpexpbf16.vhdl:314:22  */
  assign n399 = x == 9'b000001100;
  /* fpexpbf16.vhdl:315:22  */
  assign n402 = x == 9'b000001101;
  /* fpexpbf16.vhdl:316:22  */
  assign n405 = x == 9'b000001110;
  /* fpexpbf16.vhdl:317:22  */
  assign n408 = x == 9'b000001111;
  /* fpexpbf16.vhdl:318:22  */
  assign n411 = x == 9'b000010000;
  /* fpexpbf16.vhdl:319:22  */
  assign n414 = x == 9'b000010001;
  /* fpexpbf16.vhdl:320:22  */
  assign n417 = x == 9'b000010010;
  /* fpexpbf16.vhdl:321:22  */
  assign n420 = x == 9'b000010011;
  /* fpexpbf16.vhdl:322:22  */
  assign n423 = x == 9'b000010100;
  /* fpexpbf16.vhdl:323:22  */
  assign n426 = x == 9'b000010101;
  /* fpexpbf16.vhdl:324:22  */
  assign n429 = x == 9'b000010110;
  /* fpexpbf16.vhdl:325:22  */
  assign n432 = x == 9'b000010111;
  /* fpexpbf16.vhdl:326:22  */
  assign n435 = x == 9'b000011000;
  /* fpexpbf16.vhdl:327:22  */
  assign n438 = x == 9'b000011001;
  /* fpexpbf16.vhdl:328:22  */
  assign n441 = x == 9'b000011010;
  /* fpexpbf16.vhdl:329:22  */
  assign n444 = x == 9'b000011011;
  /* fpexpbf16.vhdl:330:22  */
  assign n447 = x == 9'b000011100;
  /* fpexpbf16.vhdl:331:22  */
  assign n450 = x == 9'b000011101;
  /* fpexpbf16.vhdl:332:22  */
  assign n453 = x == 9'b000011110;
  /* fpexpbf16.vhdl:333:22  */
  assign n456 = x == 9'b000011111;
  /* fpexpbf16.vhdl:334:22  */
  assign n459 = x == 9'b000100000;
  /* fpexpbf16.vhdl:335:22  */
  assign n462 = x == 9'b000100001;
  /* fpexpbf16.vhdl:336:22  */
  assign n465 = x == 9'b000100010;
  /* fpexpbf16.vhdl:337:22  */
  assign n468 = x == 9'b000100011;
  /* fpexpbf16.vhdl:338:22  */
  assign n471 = x == 9'b000100100;
  /* fpexpbf16.vhdl:339:22  */
  assign n474 = x == 9'b000100101;
  /* fpexpbf16.vhdl:340:22  */
  assign n477 = x == 9'b000100110;
  /* fpexpbf16.vhdl:341:22  */
  assign n480 = x == 9'b000100111;
  /* fpexpbf16.vhdl:342:22  */
  assign n483 = x == 9'b000101000;
  /* fpexpbf16.vhdl:343:22  */
  assign n486 = x == 9'b000101001;
  /* fpexpbf16.vhdl:344:22  */
  assign n489 = x == 9'b000101010;
  /* fpexpbf16.vhdl:345:22  */
  assign n492 = x == 9'b000101011;
  /* fpexpbf16.vhdl:346:22  */
  assign n495 = x == 9'b000101100;
  /* fpexpbf16.vhdl:347:22  */
  assign n498 = x == 9'b000101101;
  /* fpexpbf16.vhdl:348:22  */
  assign n501 = x == 9'b000101110;
  /* fpexpbf16.vhdl:349:22  */
  assign n504 = x == 9'b000101111;
  /* fpexpbf16.vhdl:350:22  */
  assign n507 = x == 9'b000110000;
  /* fpexpbf16.vhdl:351:22  */
  assign n510 = x == 9'b000110001;
  /* fpexpbf16.vhdl:352:22  */
  assign n513 = x == 9'b000110010;
  /* fpexpbf16.vhdl:353:22  */
  assign n516 = x == 9'b000110011;
  /* fpexpbf16.vhdl:354:22  */
  assign n519 = x == 9'b000110100;
  /* fpexpbf16.vhdl:355:22  */
  assign n522 = x == 9'b000110101;
  /* fpexpbf16.vhdl:356:22  */
  assign n525 = x == 9'b000110110;
  /* fpexpbf16.vhdl:357:22  */
  assign n528 = x == 9'b000110111;
  /* fpexpbf16.vhdl:358:22  */
  assign n531 = x == 9'b000111000;
  /* fpexpbf16.vhdl:359:22  */
  assign n534 = x == 9'b000111001;
  /* fpexpbf16.vhdl:360:22  */
  assign n537 = x == 9'b000111010;
  /* fpexpbf16.vhdl:361:22  */
  assign n540 = x == 9'b000111011;
  /* fpexpbf16.vhdl:362:22  */
  assign n543 = x == 9'b000111100;
  /* fpexpbf16.vhdl:363:22  */
  assign n546 = x == 9'b000111101;
  /* fpexpbf16.vhdl:364:22  */
  assign n549 = x == 9'b000111110;
  /* fpexpbf16.vhdl:365:22  */
  assign n552 = x == 9'b000111111;
  /* fpexpbf16.vhdl:366:22  */
  assign n555 = x == 9'b001000000;
  /* fpexpbf16.vhdl:367:22  */
  assign n558 = x == 9'b001000001;
  /* fpexpbf16.vhdl:368:22  */
  assign n561 = x == 9'b001000010;
  /* fpexpbf16.vhdl:369:22  */
  assign n564 = x == 9'b001000011;
  /* fpexpbf16.vhdl:370:22  */
  assign n567 = x == 9'b001000100;
  /* fpexpbf16.vhdl:371:22  */
  assign n570 = x == 9'b001000101;
  /* fpexpbf16.vhdl:372:22  */
  assign n573 = x == 9'b001000110;
  /* fpexpbf16.vhdl:373:22  */
  assign n576 = x == 9'b001000111;
  /* fpexpbf16.vhdl:374:22  */
  assign n579 = x == 9'b001001000;
  /* fpexpbf16.vhdl:375:22  */
  assign n582 = x == 9'b001001001;
  /* fpexpbf16.vhdl:376:22  */
  assign n585 = x == 9'b001001010;
  /* fpexpbf16.vhdl:377:22  */
  assign n588 = x == 9'b001001011;
  /* fpexpbf16.vhdl:378:22  */
  assign n591 = x == 9'b001001100;
  /* fpexpbf16.vhdl:379:22  */
  assign n594 = x == 9'b001001101;
  /* fpexpbf16.vhdl:380:22  */
  assign n597 = x == 9'b001001110;
  /* fpexpbf16.vhdl:381:22  */
  assign n600 = x == 9'b001001111;
  /* fpexpbf16.vhdl:382:22  */
  assign n603 = x == 9'b001010000;
  /* fpexpbf16.vhdl:383:22  */
  assign n606 = x == 9'b001010001;
  /* fpexpbf16.vhdl:384:22  */
  assign n609 = x == 9'b001010010;
  /* fpexpbf16.vhdl:385:22  */
  assign n612 = x == 9'b001010011;
  /* fpexpbf16.vhdl:386:22  */
  assign n615 = x == 9'b001010100;
  /* fpexpbf16.vhdl:387:22  */
  assign n618 = x == 9'b001010101;
  /* fpexpbf16.vhdl:388:22  */
  assign n621 = x == 9'b001010110;
  /* fpexpbf16.vhdl:389:22  */
  assign n624 = x == 9'b001010111;
  /* fpexpbf16.vhdl:390:22  */
  assign n627 = x == 9'b001011000;
  /* fpexpbf16.vhdl:391:22  */
  assign n630 = x == 9'b001011001;
  /* fpexpbf16.vhdl:392:22  */
  assign n633 = x == 9'b001011010;
  /* fpexpbf16.vhdl:393:22  */
  assign n636 = x == 9'b001011011;
  /* fpexpbf16.vhdl:394:22  */
  assign n639 = x == 9'b001011100;
  /* fpexpbf16.vhdl:395:22  */
  assign n642 = x == 9'b001011101;
  /* fpexpbf16.vhdl:396:22  */
  assign n645 = x == 9'b001011110;
  /* fpexpbf16.vhdl:397:22  */
  assign n648 = x == 9'b001011111;
  /* fpexpbf16.vhdl:398:22  */
  assign n651 = x == 9'b001100000;
  /* fpexpbf16.vhdl:399:22  */
  assign n654 = x == 9'b001100001;
  /* fpexpbf16.vhdl:400:22  */
  assign n657 = x == 9'b001100010;
  /* fpexpbf16.vhdl:401:22  */
  assign n660 = x == 9'b001100011;
  /* fpexpbf16.vhdl:402:22  */
  assign n663 = x == 9'b001100100;
  /* fpexpbf16.vhdl:403:22  */
  assign n666 = x == 9'b001100101;
  /* fpexpbf16.vhdl:404:22  */
  assign n669 = x == 9'b001100110;
  /* fpexpbf16.vhdl:405:22  */
  assign n672 = x == 9'b001100111;
  /* fpexpbf16.vhdl:406:22  */
  assign n675 = x == 9'b001101000;
  /* fpexpbf16.vhdl:407:22  */
  assign n678 = x == 9'b001101001;
  /* fpexpbf16.vhdl:408:22  */
  assign n681 = x == 9'b001101010;
  /* fpexpbf16.vhdl:409:22  */
  assign n684 = x == 9'b001101011;
  /* fpexpbf16.vhdl:410:22  */
  assign n687 = x == 9'b001101100;
  /* fpexpbf16.vhdl:411:22  */
  assign n690 = x == 9'b001101101;
  /* fpexpbf16.vhdl:412:22  */
  assign n693 = x == 9'b001101110;
  /* fpexpbf16.vhdl:413:22  */
  assign n696 = x == 9'b001101111;
  /* fpexpbf16.vhdl:414:22  */
  assign n699 = x == 9'b001110000;
  /* fpexpbf16.vhdl:415:22  */
  assign n702 = x == 9'b001110001;
  /* fpexpbf16.vhdl:416:22  */
  assign n705 = x == 9'b001110010;
  /* fpexpbf16.vhdl:417:22  */
  assign n708 = x == 9'b001110011;
  /* fpexpbf16.vhdl:418:22  */
  assign n711 = x == 9'b001110100;
  /* fpexpbf16.vhdl:419:22  */
  assign n714 = x == 9'b001110101;
  /* fpexpbf16.vhdl:420:22  */
  assign n717 = x == 9'b001110110;
  /* fpexpbf16.vhdl:421:22  */
  assign n720 = x == 9'b001110111;
  /* fpexpbf16.vhdl:422:22  */
  assign n723 = x == 9'b001111000;
  /* fpexpbf16.vhdl:423:22  */
  assign n726 = x == 9'b001111001;
  /* fpexpbf16.vhdl:424:22  */
  assign n729 = x == 9'b001111010;
  /* fpexpbf16.vhdl:425:22  */
  assign n732 = x == 9'b001111011;
  /* fpexpbf16.vhdl:426:22  */
  assign n735 = x == 9'b001111100;
  /* fpexpbf16.vhdl:427:22  */
  assign n738 = x == 9'b001111101;
  /* fpexpbf16.vhdl:428:22  */
  assign n741 = x == 9'b001111110;
  /* fpexpbf16.vhdl:429:22  */
  assign n744 = x == 9'b001111111;
  /* fpexpbf16.vhdl:430:22  */
  assign n747 = x == 9'b010000000;
  /* fpexpbf16.vhdl:431:22  */
  assign n750 = x == 9'b010000001;
  /* fpexpbf16.vhdl:432:22  */
  assign n753 = x == 9'b010000010;
  /* fpexpbf16.vhdl:433:22  */
  assign n756 = x == 9'b010000011;
  /* fpexpbf16.vhdl:434:22  */
  assign n759 = x == 9'b010000100;
  /* fpexpbf16.vhdl:435:22  */
  assign n762 = x == 9'b010000101;
  /* fpexpbf16.vhdl:436:22  */
  assign n765 = x == 9'b010000110;
  /* fpexpbf16.vhdl:437:22  */
  assign n768 = x == 9'b010000111;
  /* fpexpbf16.vhdl:438:22  */
  assign n771 = x == 9'b010001000;
  /* fpexpbf16.vhdl:439:22  */
  assign n774 = x == 9'b010001001;
  /* fpexpbf16.vhdl:440:22  */
  assign n777 = x == 9'b010001010;
  /* fpexpbf16.vhdl:441:22  */
  assign n780 = x == 9'b010001011;
  /* fpexpbf16.vhdl:442:22  */
  assign n783 = x == 9'b010001100;
  /* fpexpbf16.vhdl:443:22  */
  assign n786 = x == 9'b010001101;
  /* fpexpbf16.vhdl:444:22  */
  assign n789 = x == 9'b010001110;
  /* fpexpbf16.vhdl:445:22  */
  assign n792 = x == 9'b010001111;
  /* fpexpbf16.vhdl:446:22  */
  assign n795 = x == 9'b010010000;
  /* fpexpbf16.vhdl:447:22  */
  assign n798 = x == 9'b010010001;
  /* fpexpbf16.vhdl:448:22  */
  assign n801 = x == 9'b010010010;
  /* fpexpbf16.vhdl:449:22  */
  assign n804 = x == 9'b010010011;
  /* fpexpbf16.vhdl:450:22  */
  assign n807 = x == 9'b010010100;
  /* fpexpbf16.vhdl:451:22  */
  assign n810 = x == 9'b010010101;
  /* fpexpbf16.vhdl:452:22  */
  assign n813 = x == 9'b010010110;
  /* fpexpbf16.vhdl:453:22  */
  assign n816 = x == 9'b010010111;
  /* fpexpbf16.vhdl:454:22  */
  assign n819 = x == 9'b010011000;
  /* fpexpbf16.vhdl:455:22  */
  assign n822 = x == 9'b010011001;
  /* fpexpbf16.vhdl:456:22  */
  assign n825 = x == 9'b010011010;
  /* fpexpbf16.vhdl:457:22  */
  assign n828 = x == 9'b010011011;
  /* fpexpbf16.vhdl:458:22  */
  assign n831 = x == 9'b010011100;
  /* fpexpbf16.vhdl:459:22  */
  assign n834 = x == 9'b010011101;
  /* fpexpbf16.vhdl:460:22  */
  assign n837 = x == 9'b010011110;
  /* fpexpbf16.vhdl:461:22  */
  assign n840 = x == 9'b010011111;
  /* fpexpbf16.vhdl:462:22  */
  assign n843 = x == 9'b010100000;
  /* fpexpbf16.vhdl:463:22  */
  assign n846 = x == 9'b010100001;
  /* fpexpbf16.vhdl:464:22  */
  assign n849 = x == 9'b010100010;
  /* fpexpbf16.vhdl:465:22  */
  assign n852 = x == 9'b010100011;
  /* fpexpbf16.vhdl:466:22  */
  assign n855 = x == 9'b010100100;
  /* fpexpbf16.vhdl:467:22  */
  assign n858 = x == 9'b010100101;
  /* fpexpbf16.vhdl:468:22  */
  assign n861 = x == 9'b010100110;
  /* fpexpbf16.vhdl:469:22  */
  assign n864 = x == 9'b010100111;
  /* fpexpbf16.vhdl:470:22  */
  assign n867 = x == 9'b010101000;
  /* fpexpbf16.vhdl:471:22  */
  assign n870 = x == 9'b010101001;
  /* fpexpbf16.vhdl:472:22  */
  assign n873 = x == 9'b010101010;
  /* fpexpbf16.vhdl:473:22  */
  assign n876 = x == 9'b010101011;
  /* fpexpbf16.vhdl:474:22  */
  assign n879 = x == 9'b010101100;
  /* fpexpbf16.vhdl:475:22  */
  assign n882 = x == 9'b010101101;
  /* fpexpbf16.vhdl:476:22  */
  assign n885 = x == 9'b010101110;
  /* fpexpbf16.vhdl:477:22  */
  assign n888 = x == 9'b010101111;
  /* fpexpbf16.vhdl:478:22  */
  assign n891 = x == 9'b010110000;
  /* fpexpbf16.vhdl:479:22  */
  assign n894 = x == 9'b010110001;
  /* fpexpbf16.vhdl:480:22  */
  assign n897 = x == 9'b010110010;
  /* fpexpbf16.vhdl:481:22  */
  assign n900 = x == 9'b010110011;
  /* fpexpbf16.vhdl:482:22  */
  assign n903 = x == 9'b010110100;
  /* fpexpbf16.vhdl:483:22  */
  assign n906 = x == 9'b010110101;
  /* fpexpbf16.vhdl:484:22  */
  assign n909 = x == 9'b010110110;
  /* fpexpbf16.vhdl:485:22  */
  assign n912 = x == 9'b010110111;
  /* fpexpbf16.vhdl:486:22  */
  assign n915 = x == 9'b010111000;
  /* fpexpbf16.vhdl:487:22  */
  assign n918 = x == 9'b010111001;
  /* fpexpbf16.vhdl:488:22  */
  assign n921 = x == 9'b010111010;
  /* fpexpbf16.vhdl:489:22  */
  assign n924 = x == 9'b010111011;
  /* fpexpbf16.vhdl:490:22  */
  assign n927 = x == 9'b010111100;
  /* fpexpbf16.vhdl:491:22  */
  assign n930 = x == 9'b010111101;
  /* fpexpbf16.vhdl:492:22  */
  assign n933 = x == 9'b010111110;
  /* fpexpbf16.vhdl:493:22  */
  assign n936 = x == 9'b010111111;
  /* fpexpbf16.vhdl:494:22  */
  assign n939 = x == 9'b011000000;
  /* fpexpbf16.vhdl:495:22  */
  assign n942 = x == 9'b011000001;
  /* fpexpbf16.vhdl:496:22  */
  assign n945 = x == 9'b011000010;
  /* fpexpbf16.vhdl:497:22  */
  assign n948 = x == 9'b011000011;
  /* fpexpbf16.vhdl:498:22  */
  assign n951 = x == 9'b011000100;
  /* fpexpbf16.vhdl:499:22  */
  assign n954 = x == 9'b011000101;
  /* fpexpbf16.vhdl:500:22  */
  assign n957 = x == 9'b011000110;
  /* fpexpbf16.vhdl:501:22  */
  assign n960 = x == 9'b011000111;
  /* fpexpbf16.vhdl:502:22  */
  assign n963 = x == 9'b011001000;
  /* fpexpbf16.vhdl:503:22  */
  assign n966 = x == 9'b011001001;
  /* fpexpbf16.vhdl:504:22  */
  assign n969 = x == 9'b011001010;
  /* fpexpbf16.vhdl:505:22  */
  assign n972 = x == 9'b011001011;
  /* fpexpbf16.vhdl:506:22  */
  assign n975 = x == 9'b011001100;
  /* fpexpbf16.vhdl:507:22  */
  assign n978 = x == 9'b011001101;
  /* fpexpbf16.vhdl:508:22  */
  assign n981 = x == 9'b011001110;
  /* fpexpbf16.vhdl:509:22  */
  assign n984 = x == 9'b011001111;
  /* fpexpbf16.vhdl:510:22  */
  assign n987 = x == 9'b011010000;
  /* fpexpbf16.vhdl:511:22  */
  assign n990 = x == 9'b011010001;
  /* fpexpbf16.vhdl:512:22  */
  assign n993 = x == 9'b011010010;
  /* fpexpbf16.vhdl:513:22  */
  assign n996 = x == 9'b011010011;
  /* fpexpbf16.vhdl:514:22  */
  assign n999 = x == 9'b011010100;
  /* fpexpbf16.vhdl:515:22  */
  assign n1002 = x == 9'b011010101;
  /* fpexpbf16.vhdl:516:22  */
  assign n1005 = x == 9'b011010110;
  /* fpexpbf16.vhdl:517:22  */
  assign n1008 = x == 9'b011010111;
  /* fpexpbf16.vhdl:518:22  */
  assign n1011 = x == 9'b011011000;
  /* fpexpbf16.vhdl:519:22  */
  assign n1014 = x == 9'b011011001;
  /* fpexpbf16.vhdl:520:22  */
  assign n1017 = x == 9'b011011010;
  /* fpexpbf16.vhdl:521:22  */
  assign n1020 = x == 9'b011011011;
  /* fpexpbf16.vhdl:522:22  */
  assign n1023 = x == 9'b011011100;
  /* fpexpbf16.vhdl:523:22  */
  assign n1026 = x == 9'b011011101;
  /* fpexpbf16.vhdl:524:22  */
  assign n1029 = x == 9'b011011110;
  /* fpexpbf16.vhdl:525:22  */
  assign n1032 = x == 9'b011011111;
  /* fpexpbf16.vhdl:526:22  */
  assign n1035 = x == 9'b011100000;
  /* fpexpbf16.vhdl:527:22  */
  assign n1038 = x == 9'b011100001;
  /* fpexpbf16.vhdl:528:22  */
  assign n1041 = x == 9'b011100010;
  /* fpexpbf16.vhdl:529:22  */
  assign n1044 = x == 9'b011100011;
  /* fpexpbf16.vhdl:530:22  */
  assign n1047 = x == 9'b011100100;
  /* fpexpbf16.vhdl:531:22  */
  assign n1050 = x == 9'b011100101;
  /* fpexpbf16.vhdl:532:22  */
  assign n1053 = x == 9'b011100110;
  /* fpexpbf16.vhdl:533:22  */
  assign n1056 = x == 9'b011100111;
  /* fpexpbf16.vhdl:534:22  */
  assign n1059 = x == 9'b011101000;
  /* fpexpbf16.vhdl:535:22  */
  assign n1062 = x == 9'b011101001;
  /* fpexpbf16.vhdl:536:22  */
  assign n1065 = x == 9'b011101010;
  /* fpexpbf16.vhdl:537:22  */
  assign n1068 = x == 9'b011101011;
  /* fpexpbf16.vhdl:538:22  */
  assign n1071 = x == 9'b011101100;
  /* fpexpbf16.vhdl:539:22  */
  assign n1074 = x == 9'b011101101;
  /* fpexpbf16.vhdl:540:22  */
  assign n1077 = x == 9'b011101110;
  /* fpexpbf16.vhdl:541:22  */
  assign n1080 = x == 9'b011101111;
  /* fpexpbf16.vhdl:542:22  */
  assign n1083 = x == 9'b011110000;
  /* fpexpbf16.vhdl:543:22  */
  assign n1086 = x == 9'b011110001;
  /* fpexpbf16.vhdl:544:22  */
  assign n1089 = x == 9'b011110010;
  /* fpexpbf16.vhdl:545:22  */
  assign n1092 = x == 9'b011110011;
  /* fpexpbf16.vhdl:546:22  */
  assign n1095 = x == 9'b011110100;
  /* fpexpbf16.vhdl:547:22  */
  assign n1098 = x == 9'b011110101;
  /* fpexpbf16.vhdl:548:22  */
  assign n1101 = x == 9'b011110110;
  /* fpexpbf16.vhdl:549:22  */
  assign n1104 = x == 9'b011110111;
  /* fpexpbf16.vhdl:550:22  */
  assign n1107 = x == 9'b011111000;
  /* fpexpbf16.vhdl:551:22  */
  assign n1110 = x == 9'b011111001;
  /* fpexpbf16.vhdl:552:22  */
  assign n1113 = x == 9'b011111010;
  /* fpexpbf16.vhdl:553:22  */
  assign n1116 = x == 9'b011111011;
  /* fpexpbf16.vhdl:554:22  */
  assign n1119 = x == 9'b011111100;
  /* fpexpbf16.vhdl:555:22  */
  assign n1122 = x == 9'b011111101;
  /* fpexpbf16.vhdl:556:22  */
  assign n1125 = x == 9'b011111110;
  /* fpexpbf16.vhdl:557:22  */
  assign n1128 = x == 9'b011111111;
  /* fpexpbf16.vhdl:558:22  */
  assign n1131 = x == 9'b100000000;
  /* fpexpbf16.vhdl:559:22  */
  assign n1134 = x == 9'b100000001;
  /* fpexpbf16.vhdl:560:22  */
  assign n1137 = x == 9'b100000010;
  /* fpexpbf16.vhdl:561:22  */
  assign n1140 = x == 9'b100000011;
  /* fpexpbf16.vhdl:562:22  */
  assign n1143 = x == 9'b100000100;
  /* fpexpbf16.vhdl:563:22  */
  assign n1146 = x == 9'b100000101;
  /* fpexpbf16.vhdl:564:22  */
  assign n1149 = x == 9'b100000110;
  /* fpexpbf16.vhdl:565:22  */
  assign n1152 = x == 9'b100000111;
  /* fpexpbf16.vhdl:566:22  */
  assign n1155 = x == 9'b100001000;
  /* fpexpbf16.vhdl:567:22  */
  assign n1158 = x == 9'b100001001;
  /* fpexpbf16.vhdl:568:22  */
  assign n1161 = x == 9'b100001010;
  /* fpexpbf16.vhdl:569:22  */
  assign n1164 = x == 9'b100001011;
  /* fpexpbf16.vhdl:570:22  */
  assign n1167 = x == 9'b100001100;
  /* fpexpbf16.vhdl:571:22  */
  assign n1170 = x == 9'b100001101;
  /* fpexpbf16.vhdl:572:22  */
  assign n1173 = x == 9'b100001110;
  /* fpexpbf16.vhdl:573:22  */
  assign n1176 = x == 9'b100001111;
  /* fpexpbf16.vhdl:574:22  */
  assign n1179 = x == 9'b100010000;
  /* fpexpbf16.vhdl:575:22  */
  assign n1182 = x == 9'b100010001;
  /* fpexpbf16.vhdl:576:22  */
  assign n1185 = x == 9'b100010010;
  /* fpexpbf16.vhdl:577:22  */
  assign n1188 = x == 9'b100010011;
  /* fpexpbf16.vhdl:578:22  */
  assign n1191 = x == 9'b100010100;
  /* fpexpbf16.vhdl:579:22  */
  assign n1194 = x == 9'b100010101;
  /* fpexpbf16.vhdl:580:22  */
  assign n1197 = x == 9'b100010110;
  /* fpexpbf16.vhdl:581:22  */
  assign n1200 = x == 9'b100010111;
  /* fpexpbf16.vhdl:582:22  */
  assign n1203 = x == 9'b100011000;
  /* fpexpbf16.vhdl:583:22  */
  assign n1206 = x == 9'b100011001;
  /* fpexpbf16.vhdl:584:22  */
  assign n1209 = x == 9'b100011010;
  /* fpexpbf16.vhdl:585:22  */
  assign n1212 = x == 9'b100011011;
  /* fpexpbf16.vhdl:586:22  */
  assign n1215 = x == 9'b100011100;
  /* fpexpbf16.vhdl:587:22  */
  assign n1218 = x == 9'b100011101;
  /* fpexpbf16.vhdl:588:22  */
  assign n1221 = x == 9'b100011110;
  /* fpexpbf16.vhdl:589:22  */
  assign n1224 = x == 9'b100011111;
  /* fpexpbf16.vhdl:590:22  */
  assign n1227 = x == 9'b100100000;
  /* fpexpbf16.vhdl:591:22  */
  assign n1230 = x == 9'b100100001;
  /* fpexpbf16.vhdl:592:22  */
  assign n1233 = x == 9'b100100010;
  /* fpexpbf16.vhdl:593:22  */
  assign n1236 = x == 9'b100100011;
  /* fpexpbf16.vhdl:594:22  */
  assign n1239 = x == 9'b100100100;
  /* fpexpbf16.vhdl:595:22  */
  assign n1242 = x == 9'b100100101;
  /* fpexpbf16.vhdl:596:22  */
  assign n1245 = x == 9'b100100110;
  /* fpexpbf16.vhdl:597:22  */
  assign n1248 = x == 9'b100100111;
  /* fpexpbf16.vhdl:598:22  */
  assign n1251 = x == 9'b100101000;
  /* fpexpbf16.vhdl:599:22  */
  assign n1254 = x == 9'b100101001;
  /* fpexpbf16.vhdl:600:22  */
  assign n1257 = x == 9'b100101010;
  /* fpexpbf16.vhdl:601:22  */
  assign n1260 = x == 9'b100101011;
  /* fpexpbf16.vhdl:602:22  */
  assign n1263 = x == 9'b100101100;
  /* fpexpbf16.vhdl:603:22  */
  assign n1266 = x == 9'b100101101;
  /* fpexpbf16.vhdl:604:22  */
  assign n1269 = x == 9'b100101110;
  /* fpexpbf16.vhdl:605:22  */
  assign n1272 = x == 9'b100101111;
  /* fpexpbf16.vhdl:606:22  */
  assign n1275 = x == 9'b100110000;
  /* fpexpbf16.vhdl:607:22  */
  assign n1278 = x == 9'b100110001;
  /* fpexpbf16.vhdl:608:22  */
  assign n1281 = x == 9'b100110010;
  /* fpexpbf16.vhdl:609:22  */
  assign n1284 = x == 9'b100110011;
  /* fpexpbf16.vhdl:610:22  */
  assign n1287 = x == 9'b100110100;
  /* fpexpbf16.vhdl:611:22  */
  assign n1290 = x == 9'b100110101;
  /* fpexpbf16.vhdl:612:22  */
  assign n1293 = x == 9'b100110110;
  /* fpexpbf16.vhdl:613:22  */
  assign n1296 = x == 9'b100110111;
  /* fpexpbf16.vhdl:614:22  */
  assign n1299 = x == 9'b100111000;
  /* fpexpbf16.vhdl:615:22  */
  assign n1302 = x == 9'b100111001;
  /* fpexpbf16.vhdl:616:22  */
  assign n1305 = x == 9'b100111010;
  /* fpexpbf16.vhdl:617:22  */
  assign n1308 = x == 9'b100111011;
  /* fpexpbf16.vhdl:618:22  */
  assign n1311 = x == 9'b100111100;
  /* fpexpbf16.vhdl:619:22  */
  assign n1314 = x == 9'b100111101;
  /* fpexpbf16.vhdl:620:22  */
  assign n1317 = x == 9'b100111110;
  /* fpexpbf16.vhdl:621:22  */
  assign n1320 = x == 9'b100111111;
  /* fpexpbf16.vhdl:622:22  */
  assign n1323 = x == 9'b101000000;
  /* fpexpbf16.vhdl:623:22  */
  assign n1326 = x == 9'b101000001;
  /* fpexpbf16.vhdl:624:22  */
  assign n1329 = x == 9'b101000010;
  /* fpexpbf16.vhdl:625:22  */
  assign n1332 = x == 9'b101000011;
  /* fpexpbf16.vhdl:626:22  */
  assign n1335 = x == 9'b101000100;
  /* fpexpbf16.vhdl:627:22  */
  assign n1338 = x == 9'b101000101;
  /* fpexpbf16.vhdl:628:22  */
  assign n1341 = x == 9'b101000110;
  /* fpexpbf16.vhdl:629:22  */
  assign n1344 = x == 9'b101000111;
  /* fpexpbf16.vhdl:630:22  */
  assign n1347 = x == 9'b101001000;
  /* fpexpbf16.vhdl:631:22  */
  assign n1350 = x == 9'b101001001;
  /* fpexpbf16.vhdl:632:22  */
  assign n1353 = x == 9'b101001010;
  /* fpexpbf16.vhdl:633:22  */
  assign n1356 = x == 9'b101001011;
  /* fpexpbf16.vhdl:634:22  */
  assign n1359 = x == 9'b101001100;
  /* fpexpbf16.vhdl:635:22  */
  assign n1362 = x == 9'b101001101;
  /* fpexpbf16.vhdl:636:22  */
  assign n1365 = x == 9'b101001110;
  /* fpexpbf16.vhdl:637:22  */
  assign n1368 = x == 9'b101001111;
  /* fpexpbf16.vhdl:638:22  */
  assign n1371 = x == 9'b101010000;
  /* fpexpbf16.vhdl:639:22  */
  assign n1374 = x == 9'b101010001;
  /* fpexpbf16.vhdl:640:22  */
  assign n1377 = x == 9'b101010010;
  /* fpexpbf16.vhdl:641:22  */
  assign n1380 = x == 9'b101010011;
  /* fpexpbf16.vhdl:642:22  */
  assign n1383 = x == 9'b101010100;
  /* fpexpbf16.vhdl:643:22  */
  assign n1386 = x == 9'b101010101;
  /* fpexpbf16.vhdl:644:22  */
  assign n1389 = x == 9'b101010110;
  /* fpexpbf16.vhdl:645:22  */
  assign n1392 = x == 9'b101010111;
  /* fpexpbf16.vhdl:646:22  */
  assign n1395 = x == 9'b101011000;
  /* fpexpbf16.vhdl:647:22  */
  assign n1398 = x == 9'b101011001;
  /* fpexpbf16.vhdl:648:22  */
  assign n1401 = x == 9'b101011010;
  /* fpexpbf16.vhdl:649:22  */
  assign n1404 = x == 9'b101011011;
  /* fpexpbf16.vhdl:650:22  */
  assign n1407 = x == 9'b101011100;
  /* fpexpbf16.vhdl:651:22  */
  assign n1410 = x == 9'b101011101;
  /* fpexpbf16.vhdl:652:22  */
  assign n1413 = x == 9'b101011110;
  /* fpexpbf16.vhdl:653:22  */
  assign n1416 = x == 9'b101011111;
  /* fpexpbf16.vhdl:654:22  */
  assign n1419 = x == 9'b101100000;
  /* fpexpbf16.vhdl:655:22  */
  assign n1422 = x == 9'b101100001;
  /* fpexpbf16.vhdl:656:22  */
  assign n1425 = x == 9'b101100010;
  /* fpexpbf16.vhdl:657:22  */
  assign n1428 = x == 9'b101100011;
  /* fpexpbf16.vhdl:658:22  */
  assign n1431 = x == 9'b101100100;
  /* fpexpbf16.vhdl:659:22  */
  assign n1434 = x == 9'b101100101;
  /* fpexpbf16.vhdl:660:22  */
  assign n1437 = x == 9'b101100110;
  /* fpexpbf16.vhdl:661:22  */
  assign n1440 = x == 9'b101100111;
  /* fpexpbf16.vhdl:662:22  */
  assign n1443 = x == 9'b101101000;
  /* fpexpbf16.vhdl:663:22  */
  assign n1446 = x == 9'b101101001;
  /* fpexpbf16.vhdl:664:22  */
  assign n1449 = x == 9'b101101010;
  /* fpexpbf16.vhdl:665:22  */
  assign n1452 = x == 9'b101101011;
  /* fpexpbf16.vhdl:666:22  */
  assign n1455 = x == 9'b101101100;
  /* fpexpbf16.vhdl:667:22  */
  assign n1458 = x == 9'b101101101;
  /* fpexpbf16.vhdl:668:22  */
  assign n1461 = x == 9'b101101110;
  /* fpexpbf16.vhdl:669:22  */
  assign n1464 = x == 9'b101101111;
  /* fpexpbf16.vhdl:670:22  */
  assign n1467 = x == 9'b101110000;
  /* fpexpbf16.vhdl:671:22  */
  assign n1470 = x == 9'b101110001;
  /* fpexpbf16.vhdl:672:22  */
  assign n1473 = x == 9'b101110010;
  /* fpexpbf16.vhdl:673:22  */
  assign n1476 = x == 9'b101110011;
  /* fpexpbf16.vhdl:674:22  */
  assign n1479 = x == 9'b101110100;
  /* fpexpbf16.vhdl:675:22  */
  assign n1482 = x == 9'b101110101;
  /* fpexpbf16.vhdl:676:22  */
  assign n1485 = x == 9'b101110110;
  /* fpexpbf16.vhdl:677:22  */
  assign n1488 = x == 9'b101110111;
  /* fpexpbf16.vhdl:678:22  */
  assign n1491 = x == 9'b101111000;
  /* fpexpbf16.vhdl:679:22  */
  assign n1494 = x == 9'b101111001;
  /* fpexpbf16.vhdl:680:22  */
  assign n1497 = x == 9'b101111010;
  /* fpexpbf16.vhdl:681:22  */
  assign n1500 = x == 9'b101111011;
  /* fpexpbf16.vhdl:682:22  */
  assign n1503 = x == 9'b101111100;
  /* fpexpbf16.vhdl:683:22  */
  assign n1506 = x == 9'b101111101;
  /* fpexpbf16.vhdl:684:22  */
  assign n1509 = x == 9'b101111110;
  /* fpexpbf16.vhdl:685:22  */
  assign n1512 = x == 9'b101111111;
  /* fpexpbf16.vhdl:686:22  */
  assign n1515 = x == 9'b110000000;
  /* fpexpbf16.vhdl:687:22  */
  assign n1518 = x == 9'b110000001;
  /* fpexpbf16.vhdl:688:22  */
  assign n1521 = x == 9'b110000010;
  /* fpexpbf16.vhdl:689:22  */
  assign n1524 = x == 9'b110000011;
  /* fpexpbf16.vhdl:690:22  */
  assign n1527 = x == 9'b110000100;
  /* fpexpbf16.vhdl:691:22  */
  assign n1530 = x == 9'b110000101;
  /* fpexpbf16.vhdl:692:22  */
  assign n1533 = x == 9'b110000110;
  /* fpexpbf16.vhdl:693:22  */
  assign n1536 = x == 9'b110000111;
  /* fpexpbf16.vhdl:694:22  */
  assign n1539 = x == 9'b110001000;
  /* fpexpbf16.vhdl:695:22  */
  assign n1542 = x == 9'b110001001;
  /* fpexpbf16.vhdl:696:22  */
  assign n1545 = x == 9'b110001010;
  /* fpexpbf16.vhdl:697:22  */
  assign n1548 = x == 9'b110001011;
  /* fpexpbf16.vhdl:698:22  */
  assign n1551 = x == 9'b110001100;
  /* fpexpbf16.vhdl:699:22  */
  assign n1554 = x == 9'b110001101;
  /* fpexpbf16.vhdl:700:22  */
  assign n1557 = x == 9'b110001110;
  /* fpexpbf16.vhdl:701:22  */
  assign n1560 = x == 9'b110001111;
  /* fpexpbf16.vhdl:702:22  */
  assign n1563 = x == 9'b110010000;
  /* fpexpbf16.vhdl:703:22  */
  assign n1566 = x == 9'b110010001;
  /* fpexpbf16.vhdl:704:22  */
  assign n1569 = x == 9'b110010010;
  /* fpexpbf16.vhdl:705:22  */
  assign n1572 = x == 9'b110010011;
  /* fpexpbf16.vhdl:706:22  */
  assign n1575 = x == 9'b110010100;
  /* fpexpbf16.vhdl:707:22  */
  assign n1578 = x == 9'b110010101;
  /* fpexpbf16.vhdl:708:22  */
  assign n1581 = x == 9'b110010110;
  /* fpexpbf16.vhdl:709:22  */
  assign n1584 = x == 9'b110010111;
  /* fpexpbf16.vhdl:710:22  */
  assign n1587 = x == 9'b110011000;
  /* fpexpbf16.vhdl:711:22  */
  assign n1590 = x == 9'b110011001;
  /* fpexpbf16.vhdl:712:22  */
  assign n1593 = x == 9'b110011010;
  /* fpexpbf16.vhdl:713:22  */
  assign n1596 = x == 9'b110011011;
  /* fpexpbf16.vhdl:714:22  */
  assign n1599 = x == 9'b110011100;
  /* fpexpbf16.vhdl:715:22  */
  assign n1602 = x == 9'b110011101;
  /* fpexpbf16.vhdl:716:22  */
  assign n1605 = x == 9'b110011110;
  /* fpexpbf16.vhdl:717:22  */
  assign n1608 = x == 9'b110011111;
  /* fpexpbf16.vhdl:718:22  */
  assign n1611 = x == 9'b110100000;
  /* fpexpbf16.vhdl:719:22  */
  assign n1614 = x == 9'b110100001;
  /* fpexpbf16.vhdl:720:22  */
  assign n1617 = x == 9'b110100010;
  /* fpexpbf16.vhdl:721:22  */
  assign n1620 = x == 9'b110100011;
  /* fpexpbf16.vhdl:722:22  */
  assign n1623 = x == 9'b110100100;
  /* fpexpbf16.vhdl:723:22  */
  assign n1626 = x == 9'b110100101;
  /* fpexpbf16.vhdl:724:22  */
  assign n1629 = x == 9'b110100110;
  /* fpexpbf16.vhdl:725:22  */
  assign n1632 = x == 9'b110100111;
  /* fpexpbf16.vhdl:726:22  */
  assign n1635 = x == 9'b110101000;
  /* fpexpbf16.vhdl:727:22  */
  assign n1638 = x == 9'b110101001;
  /* fpexpbf16.vhdl:728:22  */
  assign n1641 = x == 9'b110101010;
  /* fpexpbf16.vhdl:729:22  */
  assign n1644 = x == 9'b110101011;
  /* fpexpbf16.vhdl:730:22  */
  assign n1647 = x == 9'b110101100;
  /* fpexpbf16.vhdl:731:22  */
  assign n1650 = x == 9'b110101101;
  /* fpexpbf16.vhdl:732:22  */
  assign n1653 = x == 9'b110101110;
  /* fpexpbf16.vhdl:733:22  */
  assign n1656 = x == 9'b110101111;
  /* fpexpbf16.vhdl:734:22  */
  assign n1659 = x == 9'b110110000;
  /* fpexpbf16.vhdl:735:22  */
  assign n1662 = x == 9'b110110001;
  /* fpexpbf16.vhdl:736:22  */
  assign n1665 = x == 9'b110110010;
  /* fpexpbf16.vhdl:737:22  */
  assign n1668 = x == 9'b110110011;
  /* fpexpbf16.vhdl:738:22  */
  assign n1671 = x == 9'b110110100;
  /* fpexpbf16.vhdl:739:22  */
  assign n1674 = x == 9'b110110101;
  /* fpexpbf16.vhdl:740:22  */
  assign n1677 = x == 9'b110110110;
  /* fpexpbf16.vhdl:741:22  */
  assign n1680 = x == 9'b110110111;
  /* fpexpbf16.vhdl:742:22  */
  assign n1683 = x == 9'b110111000;
  /* fpexpbf16.vhdl:743:22  */
  assign n1686 = x == 9'b110111001;
  /* fpexpbf16.vhdl:744:22  */
  assign n1689 = x == 9'b110111010;
  /* fpexpbf16.vhdl:745:22  */
  assign n1692 = x == 9'b110111011;
  /* fpexpbf16.vhdl:746:22  */
  assign n1695 = x == 9'b110111100;
  /* fpexpbf16.vhdl:747:22  */
  assign n1698 = x == 9'b110111101;
  /* fpexpbf16.vhdl:748:22  */
  assign n1701 = x == 9'b110111110;
  /* fpexpbf16.vhdl:749:22  */
  assign n1704 = x == 9'b110111111;
  /* fpexpbf16.vhdl:750:22  */
  assign n1707 = x == 9'b111000000;
  /* fpexpbf16.vhdl:751:22  */
  assign n1710 = x == 9'b111000001;
  /* fpexpbf16.vhdl:752:22  */
  assign n1713 = x == 9'b111000010;
  /* fpexpbf16.vhdl:753:22  */
  assign n1716 = x == 9'b111000011;
  /* fpexpbf16.vhdl:754:22  */
  assign n1719 = x == 9'b111000100;
  /* fpexpbf16.vhdl:755:22  */
  assign n1722 = x == 9'b111000101;
  /* fpexpbf16.vhdl:756:22  */
  assign n1725 = x == 9'b111000110;
  /* fpexpbf16.vhdl:757:22  */
  assign n1728 = x == 9'b111000111;
  /* fpexpbf16.vhdl:758:22  */
  assign n1731 = x == 9'b111001000;
  /* fpexpbf16.vhdl:759:22  */
  assign n1734 = x == 9'b111001001;
  /* fpexpbf16.vhdl:760:22  */
  assign n1737 = x == 9'b111001010;
  /* fpexpbf16.vhdl:761:22  */
  assign n1740 = x == 9'b111001011;
  /* fpexpbf16.vhdl:762:22  */
  assign n1743 = x == 9'b111001100;
  /* fpexpbf16.vhdl:763:22  */
  assign n1746 = x == 9'b111001101;
  /* fpexpbf16.vhdl:764:22  */
  assign n1749 = x == 9'b111001110;
  /* fpexpbf16.vhdl:765:22  */
  assign n1752 = x == 9'b111001111;
  /* fpexpbf16.vhdl:766:22  */
  assign n1755 = x == 9'b111010000;
  /* fpexpbf16.vhdl:767:22  */
  assign n1758 = x == 9'b111010001;
  /* fpexpbf16.vhdl:768:22  */
  assign n1761 = x == 9'b111010010;
  /* fpexpbf16.vhdl:769:22  */
  assign n1764 = x == 9'b111010011;
  /* fpexpbf16.vhdl:770:22  */
  assign n1767 = x == 9'b111010100;
  /* fpexpbf16.vhdl:771:22  */
  assign n1770 = x == 9'b111010101;
  /* fpexpbf16.vhdl:772:22  */
  assign n1773 = x == 9'b111010110;
  /* fpexpbf16.vhdl:773:22  */
  assign n1776 = x == 9'b111010111;
  /* fpexpbf16.vhdl:774:22  */
  assign n1779 = x == 9'b111011000;
  /* fpexpbf16.vhdl:775:22  */
  assign n1782 = x == 9'b111011001;
  /* fpexpbf16.vhdl:776:22  */
  assign n1785 = x == 9'b111011010;
  /* fpexpbf16.vhdl:777:22  */
  assign n1788 = x == 9'b111011011;
  /* fpexpbf16.vhdl:778:22  */
  assign n1791 = x == 9'b111011100;
  /* fpexpbf16.vhdl:779:22  */
  assign n1794 = x == 9'b111011101;
  /* fpexpbf16.vhdl:780:22  */
  assign n1797 = x == 9'b111011110;
  /* fpexpbf16.vhdl:781:22  */
  assign n1800 = x == 9'b111011111;
  /* fpexpbf16.vhdl:782:22  */
  assign n1803 = x == 9'b111100000;
  /* fpexpbf16.vhdl:783:22  */
  assign n1806 = x == 9'b111100001;
  /* fpexpbf16.vhdl:784:22  */
  assign n1809 = x == 9'b111100010;
  /* fpexpbf16.vhdl:785:22  */
  assign n1812 = x == 9'b111100011;
  /* fpexpbf16.vhdl:786:22  */
  assign n1815 = x == 9'b111100100;
  /* fpexpbf16.vhdl:787:22  */
  assign n1818 = x == 9'b111100101;
  /* fpexpbf16.vhdl:788:22  */
  assign n1821 = x == 9'b111100110;
  /* fpexpbf16.vhdl:789:22  */
  assign n1824 = x == 9'b111100111;
  /* fpexpbf16.vhdl:790:22  */
  assign n1827 = x == 9'b111101000;
  /* fpexpbf16.vhdl:791:22  */
  assign n1830 = x == 9'b111101001;
  /* fpexpbf16.vhdl:792:22  */
  assign n1833 = x == 9'b111101010;
  /* fpexpbf16.vhdl:793:22  */
  assign n1836 = x == 9'b111101011;
  /* fpexpbf16.vhdl:794:22  */
  assign n1839 = x == 9'b111101100;
  /* fpexpbf16.vhdl:795:22  */
  assign n1842 = x == 9'b111101101;
  /* fpexpbf16.vhdl:796:22  */
  assign n1845 = x == 9'b111101110;
  /* fpexpbf16.vhdl:797:22  */
  assign n1848 = x == 9'b111101111;
  /* fpexpbf16.vhdl:798:22  */
  assign n1851 = x == 9'b111110000;
  /* fpexpbf16.vhdl:799:22  */
  assign n1854 = x == 9'b111110001;
  /* fpexpbf16.vhdl:800:22  */
  assign n1857 = x == 9'b111110010;
  /* fpexpbf16.vhdl:801:22  */
  assign n1860 = x == 9'b111110011;
  /* fpexpbf16.vhdl:802:22  */
  assign n1863 = x == 9'b111110100;
  /* fpexpbf16.vhdl:803:22  */
  assign n1866 = x == 9'b111110101;
  /* fpexpbf16.vhdl:804:22  */
  assign n1869 = x == 9'b111110110;
  /* fpexpbf16.vhdl:805:22  */
  assign n1872 = x == 9'b111110111;
  /* fpexpbf16.vhdl:806:22  */
  assign n1875 = x == 9'b111111000;
  /* fpexpbf16.vhdl:807:22  */
  assign n1878 = x == 9'b111111001;
  /* fpexpbf16.vhdl:808:22  */
  assign n1881 = x == 9'b111111010;
  /* fpexpbf16.vhdl:809:22  */
  assign n1884 = x == 9'b111111011;
  /* fpexpbf16.vhdl:810:22  */
  assign n1887 = x == 9'b111111100;
  /* fpexpbf16.vhdl:811:22  */
  assign n1890 = x == 9'b111111101;
  /* fpexpbf16.vhdl:812:22  */
  assign n1893 = x == 9'b111111110;
  /* fpexpbf16.vhdl:813:22  */
  assign n1896 = x == 9'b111111111;
  assign n1898 = {n1896, n1893, n1890, n1887, n1884, n1881, n1878, n1875, n1872, n1869, n1866, n1863, n1860, n1857, n1854, n1851, n1848, n1845, n1842, n1839, n1836, n1833, n1830, n1827, n1824, n1821, n1818, n1815, n1812, n1809, n1806, n1803, n1800, n1797, n1794, n1791, n1788, n1785, n1782, n1779, n1776, n1773, n1770, n1767, n1764, n1761, n1758, n1755, n1752, n1749, n1746, n1743, n1740, n1737, n1734, n1731, n1728, n1725, n1722, n1719, n1716, n1713, n1710, n1707, n1704, n1701, n1698, n1695, n1692, n1689, n1686, n1683, n1680, n1677, n1674, n1671, n1668, n1665, n1662, n1659, n1656, n1653, n1650, n1647, n1644, n1641, n1638, n1635, n1632, n1629, n1626, n1623, n1620, n1617, n1614, n1611, n1608, n1605, n1602, n1599, n1596, n1593, n1590, n1587, n1584, n1581, n1578, n1575, n1572, n1569, n1566, n1563, n1560, n1557, n1554, n1551, n1548, n1545, n1542, n1539, n1536, n1533, n1530, n1527, n1524, n1521, n1518, n1515, n1512, n1509, n1506, n1503, n1500, n1497, n1494, n1491, n1488, n1485, n1482, n1479, n1476, n1473, n1470, n1467, n1464, n1461, n1458, n1455, n1452, n1449, n1446, n1443, n1440, n1437, n1434, n1431, n1428, n1425, n1422, n1419, n1416, n1413, n1410, n1407, n1404, n1401, n1398, n1395, n1392, n1389, n1386, n1383, n1380, n1377, n1374, n1371, n1368, n1365, n1362, n1359, n1356, n1353, n1350, n1347, n1344, n1341, n1338, n1335, n1332, n1329, n1326, n1323, n1320, n1317, n1314, n1311, n1308, n1305, n1302, n1299, n1296, n1293, n1290, n1287, n1284, n1281, n1278, n1275, n1272, n1269, n1266, n1263, n1260, n1257, n1254, n1251, n1248, n1245, n1242, n1239, n1236, n1233, n1230, n1227, n1224, n1221, n1218, n1215, n1212, n1209, n1206, n1203, n1200, n1197, n1194, n1191, n1188, n1185, n1182, n1179, n1176, n1173, n1170, n1167, n1164, n1161, n1158, n1155, n1152, n1149, n1146, n1143, n1140, n1137, n1134, n1131, n1128, n1125, n1122, n1119, n1116, n1113, n1110, n1107, n1104, n1101, n1098, n1095, n1092, n1089, n1086, n1083, n1080, n1077, n1074, n1071, n1068, n1065, n1062, n1059, n1056, n1053, n1050, n1047, n1044, n1041, n1038, n1035, n1032, n1029, n1026, n1023, n1020, n1017, n1014, n1011, n1008, n1005, n1002, n999, n996, n993, n990, n987, n984, n981, n978, n975, n972, n969, n966, n963, n960, n957, n954, n951, n948, n945, n942, n939, n936, n933, n930, n927, n924, n921, n918, n915, n912, n909, n906, n903, n900, n897, n894, n891, n888, n885, n882, n879, n876, n873, n870, n867, n864, n861, n858, n855, n852, n849, n846, n843, n840, n837, n834, n831, n828, n825, n822, n819, n816, n813, n810, n807, n804, n801, n798, n795, n792, n789, n786, n783, n780, n777, n774, n771, n768, n765, n762, n759, n756, n753, n750, n747, n744, n741, n738, n735, n732, n729, n726, n723, n720, n717, n714, n711, n708, n705, n702, n699, n696, n693, n690, n687, n684, n681, n678, n675, n672, n669, n666, n663, n660, n657, n654, n651, n648, n645, n642, n639, n636, n633, n630, n627, n624, n621, n618, n615, n612, n609, n606, n603, n600, n597, n594, n591, n588, n585, n582, n579, n576, n573, n570, n567, n564, n561, n558, n555, n552, n549, n546, n543, n540, n537, n534, n531, n528, n525, n522, n519, n516, n513, n510, n507, n504, n501, n498, n495, n492, n489, n486, n483, n480, n477, n474, n471, n468, n465, n462, n459, n456, n453, n450, n447, n444, n441, n438, n435, n432, n429, n426, n423, n420, n417, n414, n411, n408, n405, n402, n399, n396, n393, n390, n387, n384, n381, n378, n375, n372, n369, n366, n363};
  /* fpexpbf16.vhdl:301:4  */
  always @*
    case (n1898)
      512'b10000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b011111111100;
      512'b01000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b011111111000;
      512'b00100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b011111110100;
      512'b00010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b011111110000;
      512'b00001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b011111101100;
      512'b00000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b011111101000;
      512'b00000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b011111100100;
      512'b00000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b011111100000;
      512'b00000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b011111011100;
      512'b00000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b011111011000;
      512'b00000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b011111010100;
      512'b00000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b011111010001;
      512'b00000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b011111001101;
      512'b00000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b011111001001;
      512'b00000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b011111000101;
      512'b00000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b011111000001;
      512'b00000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b011110111101;
      512'b00000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b011110111001;
      512'b00000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b011110110101;
      512'b00000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b011110110010;
      512'b00000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b011110101110;
      512'b00000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b011110101010;
      512'b00000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b011110100110;
      512'b00000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b011110100010;
      512'b00000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b011110011110;
      512'b00000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b011110011011;
      512'b00000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b011110010111;
      512'b00000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b011110010011;
      512'b00000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b011110001111;
      512'b00000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b011110001011;
      512'b00000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b011110001000;
      512'b00000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b011110000100;
      512'b00000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b011110000000;
      512'b00000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b011101111100;
      512'b00000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b011101111001;
      512'b00000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b011101110101;
      512'b00000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b011101110001;
      512'b00000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b011101101110;
      512'b00000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b011101101010;
      512'b00000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b011101100110;
      512'b00000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b011101100010;
      512'b00000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b011101011111;
      512'b00000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b011101011011;
      512'b00000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b011101010111;
      512'b00000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b011101010100;
      512'b00000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b011101010000;
      512'b00000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b011101001100;
      512'b00000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b011101001001;
      512'b00000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b011101000101;
      512'b00000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b011101000001;
      512'b00000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b011100111110;
      512'b00000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b011100111010;
      512'b00000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b011100110111;
      512'b00000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b011100110011;
      512'b00000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b011100101111;
      512'b00000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b011100101100;
      512'b00000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b011100101000;
      512'b00000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b011100100101;
      512'b00000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b011100100001;
      512'b00000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b011100011110;
      512'b00000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b011100011010;
      512'b00000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b011100010110;
      512'b00000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b011100010011;
      512'b00000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b011100001111;
      512'b00000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b011100001100;
      512'b00000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b011100001000;
      512'b00000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b011100000101;
      512'b00000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b011100000001;
      512'b00000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b011011111110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b011011111010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b011011110111;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b011011110011;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b011011110000;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b011011101100;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b011011101001;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b011011100101;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b011011100010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b011011011111;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b011011011011;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b011011011000;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b011011010100;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b011011010001;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b011011001110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b011011001010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b011011000111;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b011011000011;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b011011000000;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b011010111101;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b011010111001;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b011010110110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b011010110011;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b011010101111;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b011010101100;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b011010101000;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b011010100101;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b011010100010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b011010011111;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b011010011011;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b011010011000;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b011010010101;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b011010010001;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b011010001110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b011010001011;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b011010001000;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b011010000100;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b011010000001;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b011001111110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b011001111011;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b011001110111;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b011001110100;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b011001110001;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b011001101110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b011001101010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b011001100111;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b011001100100;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b011001100001;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b011001011110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b011001011010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b011001010111;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b011001010100;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b011001010001;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b011001001110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b011001001011;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b011001000111;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b011001000100;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b011001000001;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b011000111110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b011000111011;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b011000111000;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b011000110101;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b011000110010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b011000101111;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b011000101011;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b011000101000;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b011000100101;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b011000100010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b011000011111;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b011000011100;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b011000011001;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b011000010110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b011000010011;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b011000010000;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b011000001101;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b011000001010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b011000000111;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b011000000100;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b011000000001;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b010111111110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b010111111011;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b010111111000;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b010111110101;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b010111110010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b010111101111;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b010111101100;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b010111101001;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b010111100110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b010111100011;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b010111100000;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b010111011101;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b010111011010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b010111010111;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b010111010101;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b010111010010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b010111001111;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b010111001100;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b010111001001;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b010111000110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b010111000011;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b010111000000;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b010110111101;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b010110111011;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b010110111000;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b010110110101;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b010110110010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b010110101111;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b010110101100;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b010110101001;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b010110100111;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b010110100100;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b010110100001;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b010110011110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b010110011011;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b010110011001;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b010110010110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b010110010011;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b010110010000;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b010110001101;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b010110001011;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b010110001000;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b010110000101;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b010110000010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b010110000000;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b010101111101;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b010101111010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b010101110111;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b010101110101;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b010101110010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b010101101111;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b010101101100;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b010101101010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b010101100111;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b010101100100;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b010101100010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b010101011111;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b010101011100;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b010101011010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b010101010111;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b010101010100;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b010101010010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b010101001111;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b010101001100;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b010101001010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b010101000111;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b010101000100;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b010101000010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b010100111111;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b010100111100;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b010100111010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b010100110111;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b010100110101;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b010100110010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b010100101111;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b010100101101;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b010100101010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b010100101000;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b010100100101;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b010100100011;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b010100100000;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b010100011101;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b010100011011;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b010100011000;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b010100010110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b010100010011;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b010100010001;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b010100001110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b010100001100;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b010100001001;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b010100000111;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b010100000100;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b010100000010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b010011111111;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b010011111101;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b010011111010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b010011111000;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b010011110101;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b010011110011;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b010011110000;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b010011101110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b010011101011;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b010011101001;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b010011100110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b010011100100;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b010011100001;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b010011011111;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b010011011101;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b010011011010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b110100101010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b110100100011;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b110100011101;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b110100010110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b110100010000;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b110100001001;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b110100000011;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b110011111100;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b110011110110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b110011101111;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b110011101001;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b110011100010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b110011011100;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b110011010110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b110011001111;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b110011001001;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b110011000010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b110010111100;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b110010110110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b110010101111;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b110010101001;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b110010100011;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b110010011100;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b110010010110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b110010010000;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b110010001001;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b110010000011;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b110001111101;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b110001110111;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b110001110000;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b110001101010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b110001100100;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b110001011110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b110001011000;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b110001010001;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b110001001011;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b110001000101;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b110000111111;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b110000111001;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b110000110011;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b110000101101;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b110000100111;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b110000100001;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b110000011011;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b110000010100;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b110000001110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b110000001000;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b110000000010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b101111111100;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b101111110110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b101111110000;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b101111101010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b101111100101;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b101111011111;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b101111011001;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b101111010011;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b101111001101;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b101111000111;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b101111000001;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b101110111011;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b101110110101;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b101110101111;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b101110101010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b101110100100;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b101110011110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b101110011000;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b101110010010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b101110001101;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b101110000111;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b101110000001;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b101101111011;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b101101110110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b101101110000;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b101101101010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b101101100100;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b101101011111;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b101101011001;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b101101010011;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b101101001110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b101101001000;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b101101000011;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b101100111101;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b101100110111;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b101100110010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b101100101100;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b101100100110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b101100100001;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b101100011011;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b101100010110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b101100010000;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b101100001011;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b101100000101;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b101100000000;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b101011111010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b101011110101;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b101011101111;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b101011101010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b101011100100;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b101011011111;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b101011011001;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b101011010100;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b101011001111;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b101011001001;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b101011000100;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b101010111111;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b101010111001;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b101010110100;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b101010101110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b101010101001;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b101010100100;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b101010011110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b101010011001;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b101010010100;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b101010001111;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b101010001001;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b101010000100;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b101001111111;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b101001111010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b101001110100;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b101001101111;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b101001101010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b101001100101;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b101001011111;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b101001011010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b101001010101;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b101001010000;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b101001001011;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b101001000110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b101001000001;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b101000111011;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b101000110110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b101000110001;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b101000101100;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b101000100111;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b101000100010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b101000011101;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b101000011000;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b101000010011;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b101000001110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b101000001001;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b101000000100;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b100111111111;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b100111111010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b100111110101;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b100111110000;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b100111101011;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b100111100110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b100111100001;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b100111011100;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b100111010111;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b100111010010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b100111001101;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b100111001000;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b100111000011;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b100110111111;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b100110111010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b100110110101;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b100110110000;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b100110101011;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b100110100110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b100110100010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b100110011101;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b100110011000;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b100110010011;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b100110001110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b100110001010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b100110000101;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b100110000000;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b100101111011;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b100101110111;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b100101110010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b100101101101;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b100101101000;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b100101100100;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b100101011111;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b100101011010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b100101010110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b100101010001;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b100101001100;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b100101001000;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b100101000011;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b100100111110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b100100111010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b100100110101;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b100100110001;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b100100101100;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b100100100111;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b100100100011;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b100100011110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b100100011010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b100100010101;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b100100010001;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b100100001100;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b100100001000;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b100100000011;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000: n1899 = 12'b100011111111;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000: n1899 = 12'b100011111010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000: n1899 = 12'b100011110110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000: n1899 = 12'b100011110001;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000: n1899 = 12'b100011101101;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000: n1899 = 12'b100011101000;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000: n1899 = 12'b100011100100;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000: n1899 = 12'b100011011111;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000: n1899 = 12'b100011011011;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000: n1899 = 12'b100011010111;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000: n1899 = 12'b100011010010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000: n1899 = 12'b100011001110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000: n1899 = 12'b100011001001;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000: n1899 = 12'b100011000101;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000: n1899 = 12'b100011000001;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000: n1899 = 12'b100010111100;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000: n1899 = 12'b100010111000;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000: n1899 = 12'b100010110011;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000: n1899 = 12'b100010101111;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000: n1899 = 12'b100010101011;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000: n1899 = 12'b100010100110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000: n1899 = 12'b100010100010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000: n1899 = 12'b100010011110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000: n1899 = 12'b100010011001;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000: n1899 = 12'b100010010101;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000: n1899 = 12'b100010010001;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000: n1899 = 12'b100010001101;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000: n1899 = 12'b100010001000;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000: n1899 = 12'b100010000100;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000: n1899 = 12'b100010000000;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000: n1899 = 12'b100001111100;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000: n1899 = 12'b100001110111;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000: n1899 = 12'b100001110011;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000: n1899 = 12'b100001101111;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000: n1899 = 12'b100001101011;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000: n1899 = 12'b100001100110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000: n1899 = 12'b100001100010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000: n1899 = 12'b100001011110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000: n1899 = 12'b100001011010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000: n1899 = 12'b100001010110;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000: n1899 = 12'b100001010010;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000: n1899 = 12'b100001001101;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000: n1899 = 12'b100001001001;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000: n1899 = 12'b100001000101;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000: n1899 = 12'b100001000001;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000: n1899 = 12'b100000111101;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000: n1899 = 12'b100000111001;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000: n1899 = 12'b100000110101;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000: n1899 = 12'b100000110001;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000: n1899 = 12'b100000101100;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000: n1899 = 12'b100000101000;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000: n1899 = 12'b100000100100;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000: n1899 = 12'b100000100000;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000: n1899 = 12'b100000011100;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000: n1899 = 12'b100000011000;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000: n1899 = 12'b100000010100;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000: n1899 = 12'b100000010000;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000: n1899 = 12'b100000001100;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100: n1899 = 12'b100000001000;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010: n1899 = 12'b100000000100;
      512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001: n1899 = 12'b100000000000;
      default: n1899 = 12'bX;
    endcase
endmodule

module intadder_9_freq500_uid33
  (input  clk,
   input  [8:0] x,
   input  [8:0] y,
   input  cin,
   output [8:0] r);
  wire cin_1;
  wire cin_1_d1;
  wire cin_1_d2;
  wire cin_1_d3;
  wire [9:0] x_1;
  wire [9:0] x_1_d1;
  wire [9:0] x_1_d2;
  wire [9:0] y_1;
  wire [9:0] s_1;
  wire [8:0] r_1;
  wire [9:0] n348;
  wire [9:0] n350;
  wire [9:0] n351;
  wire [9:0] n352;
  wire [9:0] n353;
  wire [8:0] n354;
  reg n355;
  reg n356;
  reg n357;
  reg [9:0] n358;
  reg [9:0] n359;
  assign r = r_1; //(module output)
  /* fpexpbf16.vhdl:1378:15  */
  assign cin_1_d1 = n355; // (signal)
  /* fpexpbf16.vhdl:1378:25  */
  assign cin_1_d2 = n356; // (signal)
  /* fpexpbf16.vhdl:1378:35  */
  assign cin_1_d3 = n357; // (signal)
  /* fpexpbf16.vhdl:1380:8  */
  assign x_1 = n348; // (signal)
  /* fpexpbf16.vhdl:1380:13  */
  assign x_1_d1 = n358; // (signal)
  /* fpexpbf16.vhdl:1380:21  */
  assign x_1_d2 = n359; // (signal)
  /* fpexpbf16.vhdl:1382:8  */
  assign y_1 = n350; // (signal)
  /* fpexpbf16.vhdl:1384:8  */
  assign s_1 = n353; // (signal)
  /* fpexpbf16.vhdl:1386:8  */
  assign r_1 = n354; // (signal)
  /* fpexpbf16.vhdl:1400:15  */
  assign n348 = {1'b0, x};
  /* fpexpbf16.vhdl:1401:15  */
  assign n350 = {1'b0, y};
  /* fpexpbf16.vhdl:1402:18  */
  assign n351 = x_1_d2 + y_1;
  /* fpexpbf16.vhdl:1402:24  */
  assign n352 = {9'b0, cin_1_d3};  //  uext
  /* fpexpbf16.vhdl:1402:24  */
  assign n353 = n351 + n352;
  /* fpexpbf16.vhdl:1403:14  */
  assign n354 = s_1[8:0]; // extract
  /* fpexpbf16.vhdl:1391:10  */
  always @(posedge clk)
    n355 <= cin_1;
  /* fpexpbf16.vhdl:1391:10  */
  always @(posedge clk)
    n356 <= cin_1_d1;
  /* fpexpbf16.vhdl:1391:10  */
  always @(posedge clk)
    n357 <= cin_1_d2;
  /* fpexpbf16.vhdl:1391:10  */
  always @(posedge clk)
    n358 <= x_1;
  /* fpexpbf16.vhdl:1391:10  */
  always @(posedge clk)
    n359 <= x_1_d1;
endmodule

module fixrealkcm_freq500_uid20
  (input  clk,
   input  [7:0] x,
   output [16:0] r);
  wire [4:0] fixrealkcm_freq500_uid20_a0;
  wire [16:0] fixrealkcm_freq500_uid20_t0;
  wire [16:0] fixrealkcm_freq500_uid20_t0_copy24;
  wire bh21_w0_0;
  wire bh21_w1_0;
  wire bh21_w2_0;
  wire bh21_w3_0;
  wire bh21_w4_0;
  wire bh21_w5_0;
  wire bh21_w6_0;
  wire bh21_w7_0;
  wire bh21_w8_0;
  wire bh21_w9_0;
  wire bh21_w10_0;
  wire bh21_w11_0;
  wire bh21_w12_0;
  wire bh21_w13_0;
  wire bh21_w14_0;
  wire bh21_w15_0;
  wire bh21_w16_0;
  wire [2:0] fixrealkcm_freq500_uid20_a1;
  wire [11:0] fixrealkcm_freq500_uid20_t1;
  wire [11:0] fixrealkcm_freq500_uid20_t1_copy27;
  wire bh21_w0_1;
  wire bh21_w1_1;
  wire bh21_w2_1;
  wire bh21_w3_1;
  wire bh21_w4_1;
  wire bh21_w5_1;
  wire bh21_w6_1;
  wire bh21_w7_1;
  wire bh21_w8_1;
  wire bh21_w9_1;
  wire bh21_w10_1;
  wire bh21_w11_1;
  wire [16:0] bitheapfinaladd_bh21_in0;
  wire [16:0] bitheapfinaladd_bh21_in1;
  wire bitheapfinaladd_bh21_cin;
  wire [16:0] bitheapfinaladd_bh21_out;
  wire [16:0] bitheapresult_bh21;
  wire [16:0] outres;
  wire [4:0] n266;
  wire [16:0] fixrealkcm_freq500_uid20_table0_n267;
  wire n270;
  wire n271;
  wire n272;
  wire n273;
  wire n274;
  wire n275;
  wire n276;
  wire n277;
  wire n278;
  wire n279;
  wire n280;
  wire n281;
  wire n282;
  wire n283;
  wire n284;
  wire n285;
  wire n286;
  wire [2:0] n287;
  wire [11:0] fixrealkcm_freq500_uid20_table1_n288;
  wire n291;
  wire n292;
  wire n293;
  wire n294;
  wire n295;
  wire n296;
  wire n297;
  wire n298;
  wire n299;
  wire n300;
  wire n301;
  wire n302;
  wire [1:0] n304;
  wire [2:0] n305;
  wire [3:0] n306;
  wire [4:0] n307;
  wire [5:0] n308;
  wire [6:0] n309;
  wire [7:0] n310;
  wire [8:0] n311;
  wire [9:0] n312;
  wire [10:0] n313;
  wire [11:0] n314;
  wire [12:0] n315;
  wire [13:0] n316;
  wire [14:0] n317;
  wire [15:0] n318;
  wire [16:0] n319;
  wire [5:0] n321;
  wire [6:0] n322;
  wire [7:0] n323;
  wire [8:0] n324;
  wire [9:0] n325;
  wire [10:0] n326;
  wire [11:0] n327;
  wire [12:0] n328;
  wire [13:0] n329;
  wire [14:0] n330;
  wire [15:0] n331;
  wire [16:0] n332;
  wire [16:0] bitheapfinaladd_bh21_n334;
  assign r = outres; //(module output)
  /* fpexpbf16.vhdl:1203:8  */
  assign fixrealkcm_freq500_uid20_a0 = n266; // (signal)
  /* fpexpbf16.vhdl:1205:8  */
  assign fixrealkcm_freq500_uid20_t0 = fixrealkcm_freq500_uid20_t0_copy24; // (signal)
  /* fpexpbf16.vhdl:1207:8  */
  assign fixrealkcm_freq500_uid20_t0_copy24 = fixrealkcm_freq500_uid20_table0_n267; // (signal)
  /* fpexpbf16.vhdl:1209:8  */
  assign bh21_w0_0 = n270; // (signal)
  /* fpexpbf16.vhdl:1211:8  */
  assign bh21_w1_0 = n271; // (signal)
  /* fpexpbf16.vhdl:1213:8  */
  assign bh21_w2_0 = n272; // (signal)
  /* fpexpbf16.vhdl:1215:8  */
  assign bh21_w3_0 = n273; // (signal)
  /* fpexpbf16.vhdl:1217:8  */
  assign bh21_w4_0 = n274; // (signal)
  /* fpexpbf16.vhdl:1219:8  */
  assign bh21_w5_0 = n275; // (signal)
  /* fpexpbf16.vhdl:1221:8  */
  assign bh21_w6_0 = n276; // (signal)
  /* fpexpbf16.vhdl:1223:8  */
  assign bh21_w7_0 = n277; // (signal)
  /* fpexpbf16.vhdl:1225:8  */
  assign bh21_w8_0 = n278; // (signal)
  /* fpexpbf16.vhdl:1227:8  */
  assign bh21_w9_0 = n279; // (signal)
  /* fpexpbf16.vhdl:1229:8  */
  assign bh21_w10_0 = n280; // (signal)
  /* fpexpbf16.vhdl:1231:8  */
  assign bh21_w11_0 = n281; // (signal)
  /* fpexpbf16.vhdl:1233:8  */
  assign bh21_w12_0 = n282; // (signal)
  /* fpexpbf16.vhdl:1235:8  */
  assign bh21_w13_0 = n283; // (signal)
  /* fpexpbf16.vhdl:1237:8  */
  assign bh21_w14_0 = n284; // (signal)
  /* fpexpbf16.vhdl:1239:8  */
  assign bh21_w15_0 = n285; // (signal)
  /* fpexpbf16.vhdl:1331:35  */
  assign bh21_w16_0 = n286; // (signal)
  /* fpexpbf16.vhdl:1243:8  */
  assign fixrealkcm_freq500_uid20_a1 = n287; // (signal)
  /* fpexpbf16.vhdl:1245:8  */
  assign fixrealkcm_freq500_uid20_t1 = fixrealkcm_freq500_uid20_t1_copy27; // (signal)
  /* fpexpbf16.vhdl:1247:8  */
  assign fixrealkcm_freq500_uid20_t1_copy27 = fixrealkcm_freq500_uid20_table1_n288; // (signal)
  /* fpexpbf16.vhdl:1249:8  */
  assign bh21_w0_1 = n291; // (signal)
  /* fpexpbf16.vhdl:1251:8  */
  assign bh21_w1_1 = n292; // (signal)
  /* fpexpbf16.vhdl:1253:8  */
  assign bh21_w2_1 = n293; // (signal)
  /* fpexpbf16.vhdl:1255:8  */
  assign bh21_w3_1 = n294; // (signal)
  /* fpexpbf16.vhdl:1257:8  */
  assign bh21_w4_1 = n295; // (signal)
  /* fpexpbf16.vhdl:1259:8  */
  assign bh21_w5_1 = n296; // (signal)
  /* fpexpbf16.vhdl:1261:8  */
  assign bh21_w6_1 = n297; // (signal)
  /* fpexpbf16.vhdl:1263:8  */
  assign bh21_w7_1 = n298; // (signal)
  /* fpexpbf16.vhdl:1265:8  */
  assign bh21_w8_1 = n299; // (signal)
  /* fpexpbf16.vhdl:1267:8  */
  assign bh21_w9_1 = n300; // (signal)
  /* fpexpbf16.vhdl:1269:8  */
  assign bh21_w10_1 = n301; // (signal)
  /* fpexpbf16.vhdl:1271:8  */
  assign bh21_w11_1 = n302; // (signal)
  /* fpexpbf16.vhdl:1273:8  */
  assign bitheapfinaladd_bh21_in0 = n319; // (signal)
  /* fpexpbf16.vhdl:1275:8  */
  assign bitheapfinaladd_bh21_in1 = n332; // (signal)
  /* fpexpbf16.vhdl:1277:8  */
  assign bitheapfinaladd_bh21_cin = 1'b0; // (signal)
  /* fpexpbf16.vhdl:1279:8  */
  assign bitheapfinaladd_bh21_out = bitheapfinaladd_bh21_n334; // (signal)
  /* fpexpbf16.vhdl:1281:8  */
  assign bitheapresult_bh21 = bitheapfinaladd_bh21_out; // (signal)
  /* fpexpbf16.vhdl:1283:8  */
  assign outres = bitheapresult_bh21; // (signal)
  /* fpexpbf16.vhdl:1287:36  */
  assign n266 = x[7:3]; // extract
  /* fpexpbf16.vhdl:1288:4  */
  fixrealkcm_freq500_uid20_t0_freq500_uid23 fixrealkcm_freq500_uid20_table0 (
    .x(fixrealkcm_freq500_uid20_a0),
    .y(fixrealkcm_freq500_uid20_table0_n267));
  /* fpexpbf16.vhdl:1292:44  */
  assign n270 = fixrealkcm_freq500_uid20_t0[0]; // extract
  /* fpexpbf16.vhdl:1293:44  */
  assign n271 = fixrealkcm_freq500_uid20_t0[1]; // extract
  /* fpexpbf16.vhdl:1294:44  */
  assign n272 = fixrealkcm_freq500_uid20_t0[2]; // extract
  /* fpexpbf16.vhdl:1295:44  */
  assign n273 = fixrealkcm_freq500_uid20_t0[3]; // extract
  /* fpexpbf16.vhdl:1296:44  */
  assign n274 = fixrealkcm_freq500_uid20_t0[4]; // extract
  /* fpexpbf16.vhdl:1297:44  */
  assign n275 = fixrealkcm_freq500_uid20_t0[5]; // extract
  /* fpexpbf16.vhdl:1298:44  */
  assign n276 = fixrealkcm_freq500_uid20_t0[6]; // extract
  /* fpexpbf16.vhdl:1299:44  */
  assign n277 = fixrealkcm_freq500_uid20_t0[7]; // extract
  /* fpexpbf16.vhdl:1300:44  */
  assign n278 = fixrealkcm_freq500_uid20_t0[8]; // extract
  /* fpexpbf16.vhdl:1301:44  */
  assign n279 = fixrealkcm_freq500_uid20_t0[9]; // extract
  /* fpexpbf16.vhdl:1302:45  */
  assign n280 = fixrealkcm_freq500_uid20_t0[10]; // extract
  /* fpexpbf16.vhdl:1303:45  */
  assign n281 = fixrealkcm_freq500_uid20_t0[11]; // extract
  /* fpexpbf16.vhdl:1304:45  */
  assign n282 = fixrealkcm_freq500_uid20_t0[12]; // extract
  /* fpexpbf16.vhdl:1305:45  */
  assign n283 = fixrealkcm_freq500_uid20_t0[13]; // extract
  /* fpexpbf16.vhdl:1306:45  */
  assign n284 = fixrealkcm_freq500_uid20_t0[14]; // extract
  /* fpexpbf16.vhdl:1307:45  */
  assign n285 = fixrealkcm_freq500_uid20_t0[15]; // extract
  /* fpexpbf16.vhdl:1308:45  */
  assign n286 = fixrealkcm_freq500_uid20_t0[16]; // extract
  /* fpexpbf16.vhdl:1309:36  */
  assign n287 = x[2:0]; // extract
  /* fpexpbf16.vhdl:1310:4  */
  fixrealkcm_freq500_uid20_t1_freq500_uid26 fixrealkcm_freq500_uid20_table1 (
    .x(fixrealkcm_freq500_uid20_a1),
    .y(fixrealkcm_freq500_uid20_table1_n288));
  /* fpexpbf16.vhdl:1314:44  */
  assign n291 = fixrealkcm_freq500_uid20_t1[0]; // extract
  /* fpexpbf16.vhdl:1315:44  */
  assign n292 = fixrealkcm_freq500_uid20_t1[1]; // extract
  /* fpexpbf16.vhdl:1316:44  */
  assign n293 = fixrealkcm_freq500_uid20_t1[2]; // extract
  /* fpexpbf16.vhdl:1317:44  */
  assign n294 = fixrealkcm_freq500_uid20_t1[3]; // extract
  /* fpexpbf16.vhdl:1318:44  */
  assign n295 = fixrealkcm_freq500_uid20_t1[4]; // extract
  /* fpexpbf16.vhdl:1319:44  */
  assign n296 = fixrealkcm_freq500_uid20_t1[5]; // extract
  /* fpexpbf16.vhdl:1320:44  */
  assign n297 = fixrealkcm_freq500_uid20_t1[6]; // extract
  /* fpexpbf16.vhdl:1321:44  */
  assign n298 = fixrealkcm_freq500_uid20_t1[7]; // extract
  /* fpexpbf16.vhdl:1322:44  */
  assign n299 = fixrealkcm_freq500_uid20_t1[8]; // extract
  /* fpexpbf16.vhdl:1323:44  */
  assign n300 = fixrealkcm_freq500_uid20_t1[9]; // extract
  /* fpexpbf16.vhdl:1324:45  */
  assign n301 = fixrealkcm_freq500_uid20_t1[10]; // extract
  /* fpexpbf16.vhdl:1325:45  */
  assign n302 = fixrealkcm_freq500_uid20_t1[11]; // extract
  /* fpexpbf16.vhdl:1331:48  */
  assign n304 = {bh21_w16_0, bh21_w15_0};
  /* fpexpbf16.vhdl:1331:61  */
  assign n305 = {n304, bh21_w14_0};
  /* fpexpbf16.vhdl:1331:74  */
  assign n306 = {n305, bh21_w13_0};
  /* fpexpbf16.vhdl:1331:87  */
  assign n307 = {n306, bh21_w12_0};
  /* fpexpbf16.vhdl:1331:100  */
  assign n308 = {n307, bh21_w11_0};
  /* fpexpbf16.vhdl:1331:113  */
  assign n309 = {n308, bh21_w10_0};
  /* fpexpbf16.vhdl:1331:126  */
  assign n310 = {n309, bh21_w9_0};
  /* fpexpbf16.vhdl:1331:138  */
  assign n311 = {n310, bh21_w8_0};
  /* fpexpbf16.vhdl:1331:150  */
  assign n312 = {n311, bh21_w7_0};
  /* fpexpbf16.vhdl:1331:162  */
  assign n313 = {n312, bh21_w6_0};
  /* fpexpbf16.vhdl:1331:174  */
  assign n314 = {n313, bh21_w5_0};
  /* fpexpbf16.vhdl:1331:186  */
  assign n315 = {n314, bh21_w4_0};
  /* fpexpbf16.vhdl:1331:198  */
  assign n316 = {n315, bh21_w3_0};
  /* fpexpbf16.vhdl:1331:210  */
  assign n317 = {n316, bh21_w2_0};
  /* fpexpbf16.vhdl:1331:222  */
  assign n318 = {n317, bh21_w1_0};
  /* fpexpbf16.vhdl:1331:234  */
  assign n319 = {n318, bh21_w0_0};
  /* fpexpbf16.vhdl:1332:60  */
  assign n321 = {5'b00000, bh21_w11_1};
  /* fpexpbf16.vhdl:1332:73  */
  assign n322 = {n321, bh21_w10_1};
  /* fpexpbf16.vhdl:1332:86  */
  assign n323 = {n322, bh21_w9_1};
  /* fpexpbf16.vhdl:1332:98  */
  assign n324 = {n323, bh21_w8_1};
  /* fpexpbf16.vhdl:1332:110  */
  assign n325 = {n324, bh21_w7_1};
  /* fpexpbf16.vhdl:1332:122  */
  assign n326 = {n325, bh21_w6_1};
  /* fpexpbf16.vhdl:1332:134  */
  assign n327 = {n326, bh21_w5_1};
  /* fpexpbf16.vhdl:1332:146  */
  assign n328 = {n327, bh21_w4_1};
  /* fpexpbf16.vhdl:1332:158  */
  assign n329 = {n328, bh21_w3_1};
  /* fpexpbf16.vhdl:1332:170  */
  assign n330 = {n329, bh21_w2_1};
  /* fpexpbf16.vhdl:1332:182  */
  assign n331 = {n330, bh21_w1_1};
  /* fpexpbf16.vhdl:1332:194  */
  assign n332 = {n331, bh21_w0_1};
  /* fpexpbf16.vhdl:1335:4  */
  intadder_17_freq500_uid30 bitheapfinaladd_bh21 (
    .clk(clk),
    .x(bitheapfinaladd_bh21_in0),
    .y(bitheapfinaladd_bh21_in1),
    .cin(bitheapfinaladd_bh21_cin),
    .r(bitheapfinaladd_bh21_n334));
endmodule

module fixrealkcm_freq500_uid8
  (input  clk,
   input  [9:0] x,
   output [7:0] r);
  wire [4:0] fixrealkcm_freq500_uid8_a0;
  wire [11:0] fixrealkcm_freq500_uid8_t0;
  wire [11:0] fixrealkcm_freq500_uid8_t0_copy12;
  wire bh9_w0_0;
  wire bh9_w1_0;
  wire bh9_w2_0;
  wire bh9_w3_0;
  wire bh9_w4_0;
  wire bh9_w5_0;
  wire bh9_w6_0;
  wire bh9_w7_0;
  wire bh9_w8_0;
  wire bh9_w9_0;
  wire bh9_w10_0;
  wire bh9_w11_0;
  wire [4:0] fixrealkcm_freq500_uid8_a1;
  wire [6:0] fixrealkcm_freq500_uid8_t1;
  wire [6:0] fixrealkcm_freq500_uid8_t1_copy15;
  wire bh9_w0_1;
  wire bh9_w1_1;
  wire bh9_w2_1;
  wire bh9_w3_1;
  wire bh9_w4_1;
  wire bh9_w5_1;
  wire bh9_w6_1;
  wire [11:0] bitheapfinaladd_bh9_in0;
  wire [11:0] bitheapfinaladd_bh9_in1;
  wire bitheapfinaladd_bh9_cin;
  wire [11:0] bitheapfinaladd_bh9_out;
  wire [11:0] bitheapresult_bh9;
  wire [11:0] outres;
  wire [4:0] n213;
  wire [11:0] fixrealkcm_freq500_uid8_table0_n214;
  wire n217;
  wire n218;
  wire n219;
  wire n220;
  wire n221;
  wire n222;
  wire n223;
  wire n224;
  wire n225;
  wire n226;
  wire n227;
  wire n228;
  wire [4:0] n229;
  wire [6:0] fixrealkcm_freq500_uid8_table1_n230;
  wire n233;
  wire n234;
  wire n235;
  wire n236;
  wire n237;
  wire n238;
  wire n239;
  wire [1:0] n241;
  wire [2:0] n242;
  wire [3:0] n243;
  wire [4:0] n244;
  wire [5:0] n245;
  wire [6:0] n246;
  wire [7:0] n247;
  wire [8:0] n248;
  wire [9:0] n249;
  wire [10:0] n250;
  wire [11:0] n251;
  wire [5:0] n253;
  wire [6:0] n254;
  wire [7:0] n255;
  wire [8:0] n256;
  wire [9:0] n257;
  wire [10:0] n258;
  wire [11:0] n259;
  wire [11:0] bitheapfinaladd_bh9_n261;
  wire [7:0] n264;
  assign r = n264; //(module output)
  /* fpexpbf16.vhdl:987:8  */
  assign fixrealkcm_freq500_uid8_a0 = n213; // (signal)
  /* fpexpbf16.vhdl:989:8  */
  assign fixrealkcm_freq500_uid8_t0 = fixrealkcm_freq500_uid8_t0_copy12; // (signal)
  /* fpexpbf16.vhdl:991:8  */
  assign fixrealkcm_freq500_uid8_t0_copy12 = fixrealkcm_freq500_uid8_table0_n214; // (signal)
  /* fpexpbf16.vhdl:993:8  */
  assign bh9_w0_0 = n217; // (signal)
  /* fpexpbf16.vhdl:995:8  */
  assign bh9_w1_0 = n218; // (signal)
  /* fpexpbf16.vhdl:997:8  */
  assign bh9_w2_0 = n219; // (signal)
  /* fpexpbf16.vhdl:999:8  */
  assign bh9_w3_0 = n220; // (signal)
  /* fpexpbf16.vhdl:1001:8  */
  assign bh9_w4_0 = n221; // (signal)
  /* fpexpbf16.vhdl:1003:8  */
  assign bh9_w5_0 = n222; // (signal)
  /* fpexpbf16.vhdl:1005:8  */
  assign bh9_w6_0 = n223; // (signal)
  /* fpexpbf16.vhdl:1007:8  */
  assign bh9_w7_0 = n224; // (signal)
  /* fpexpbf16.vhdl:1009:8  */
  assign bh9_w8_0 = n225; // (signal)
  /* fpexpbf16.vhdl:1011:8  */
  assign bh9_w9_0 = n226; // (signal)
  /* fpexpbf16.vhdl:1013:8  */
  assign bh9_w10_0 = n227; // (signal)
  /* fpexpbf16.vhdl:1085:34  */
  assign bh9_w11_0 = n228; // (signal)
  /* fpexpbf16.vhdl:1017:8  */
  assign fixrealkcm_freq500_uid8_a1 = n229; // (signal)
  /* fpexpbf16.vhdl:1019:8  */
  assign fixrealkcm_freq500_uid8_t1 = fixrealkcm_freq500_uid8_t1_copy15; // (signal)
  /* fpexpbf16.vhdl:1021:8  */
  assign fixrealkcm_freq500_uid8_t1_copy15 = fixrealkcm_freq500_uid8_table1_n230; // (signal)
  /* fpexpbf16.vhdl:1023:8  */
  assign bh9_w0_1 = n233; // (signal)
  /* fpexpbf16.vhdl:1025:8  */
  assign bh9_w1_1 = n234; // (signal)
  /* fpexpbf16.vhdl:1027:8  */
  assign bh9_w2_1 = n235; // (signal)
  /* fpexpbf16.vhdl:1029:8  */
  assign bh9_w3_1 = n236; // (signal)
  /* fpexpbf16.vhdl:1031:8  */
  assign bh9_w4_1 = n237; // (signal)
  /* fpexpbf16.vhdl:1033:8  */
  assign bh9_w5_1 = n238; // (signal)
  /* fpexpbf16.vhdl:1035:8  */
  assign bh9_w6_1 = n239; // (signal)
  /* fpexpbf16.vhdl:1037:8  */
  assign bitheapfinaladd_bh9_in0 = n251; // (signal)
  /* fpexpbf16.vhdl:1039:8  */
  assign bitheapfinaladd_bh9_in1 = n259; // (signal)
  /* fpexpbf16.vhdl:1041:8  */
  assign bitheapfinaladd_bh9_cin = 1'b0; // (signal)
  /* fpexpbf16.vhdl:1043:8  */
  assign bitheapfinaladd_bh9_out = bitheapfinaladd_bh9_n261; // (signal)
  /* fpexpbf16.vhdl:1045:8  */
  assign bitheapresult_bh9 = bitheapfinaladd_bh9_out; // (signal)
  /* fpexpbf16.vhdl:1047:8  */
  assign outres = bitheapresult_bh9; // (signal)
  /* fpexpbf16.vhdl:1051:35  */
  assign n213 = x[9:5]; // extract
  /* fpexpbf16.vhdl:1052:4  */
  fixrealkcm_freq500_uid8_t0_freq500_uid11 fixrealkcm_freq500_uid8_table0 (
    .x(fixrealkcm_freq500_uid8_a0),
    .y(fixrealkcm_freq500_uid8_table0_n214));
  /* fpexpbf16.vhdl:1056:42  */
  assign n217 = fixrealkcm_freq500_uid8_t0[0]; // extract
  /* fpexpbf16.vhdl:1057:42  */
  assign n218 = fixrealkcm_freq500_uid8_t0[1]; // extract
  /* fpexpbf16.vhdl:1058:42  */
  assign n219 = fixrealkcm_freq500_uid8_t0[2]; // extract
  /* fpexpbf16.vhdl:1059:42  */
  assign n220 = fixrealkcm_freq500_uid8_t0[3]; // extract
  /* fpexpbf16.vhdl:1060:42  */
  assign n221 = fixrealkcm_freq500_uid8_t0[4]; // extract
  /* fpexpbf16.vhdl:1061:42  */
  assign n222 = fixrealkcm_freq500_uid8_t0[5]; // extract
  /* fpexpbf16.vhdl:1062:42  */
  assign n223 = fixrealkcm_freq500_uid8_t0[6]; // extract
  /* fpexpbf16.vhdl:1063:42  */
  assign n224 = fixrealkcm_freq500_uid8_t0[7]; // extract
  /* fpexpbf16.vhdl:1064:42  */
  assign n225 = fixrealkcm_freq500_uid8_t0[8]; // extract
  /* fpexpbf16.vhdl:1065:42  */
  assign n226 = fixrealkcm_freq500_uid8_t0[9]; // extract
  /* fpexpbf16.vhdl:1066:43  */
  assign n227 = fixrealkcm_freq500_uid8_t0[10]; // extract
  /* fpexpbf16.vhdl:1067:43  */
  assign n228 = fixrealkcm_freq500_uid8_t0[11]; // extract
  /* fpexpbf16.vhdl:1068:35  */
  assign n229 = x[4:0]; // extract
  /* fpexpbf16.vhdl:1069:4  */
  fixrealkcm_freq500_uid8_t1_freq500_uid14 fixrealkcm_freq500_uid8_table1 (
    .x(fixrealkcm_freq500_uid8_a1),
    .y(fixrealkcm_freq500_uid8_table1_n230));
  /* fpexpbf16.vhdl:1073:42  */
  assign n233 = fixrealkcm_freq500_uid8_t1[0]; // extract
  /* fpexpbf16.vhdl:1074:42  */
  assign n234 = fixrealkcm_freq500_uid8_t1[1]; // extract
  /* fpexpbf16.vhdl:1075:42  */
  assign n235 = fixrealkcm_freq500_uid8_t1[2]; // extract
  /* fpexpbf16.vhdl:1076:42  */
  assign n236 = fixrealkcm_freq500_uid8_t1[3]; // extract
  /* fpexpbf16.vhdl:1077:42  */
  assign n237 = fixrealkcm_freq500_uid8_t1[4]; // extract
  /* fpexpbf16.vhdl:1078:42  */
  assign n238 = fixrealkcm_freq500_uid8_t1[5]; // extract
  /* fpexpbf16.vhdl:1079:42  */
  assign n239 = fixrealkcm_freq500_uid8_t1[6]; // extract
  /* fpexpbf16.vhdl:1085:46  */
  assign n241 = {bh9_w11_0, bh9_w10_0};
  /* fpexpbf16.vhdl:1085:58  */
  assign n242 = {n241, bh9_w9_0};
  /* fpexpbf16.vhdl:1085:69  */
  assign n243 = {n242, bh9_w8_0};
  /* fpexpbf16.vhdl:1085:80  */
  assign n244 = {n243, bh9_w7_0};
  /* fpexpbf16.vhdl:1085:91  */
  assign n245 = {n244, bh9_w6_1};
  /* fpexpbf16.vhdl:1085:102  */
  assign n246 = {n245, bh9_w5_1};
  /* fpexpbf16.vhdl:1085:113  */
  assign n247 = {n246, bh9_w4_1};
  /* fpexpbf16.vhdl:1085:124  */
  assign n248 = {n247, bh9_w3_1};
  /* fpexpbf16.vhdl:1085:135  */
  assign n249 = {n248, bh9_w2_1};
  /* fpexpbf16.vhdl:1085:146  */
  assign n250 = {n249, bh9_w1_1};
  /* fpexpbf16.vhdl:1085:157  */
  assign n251 = {n250, bh9_w0_1};
  /* fpexpbf16.vhdl:1086:59  */
  assign n253 = {5'b00000, bh9_w6_0};
  /* fpexpbf16.vhdl:1086:70  */
  assign n254 = {n253, bh9_w5_0};
  /* fpexpbf16.vhdl:1086:81  */
  assign n255 = {n254, bh9_w4_0};
  /* fpexpbf16.vhdl:1086:92  */
  assign n256 = {n255, bh9_w3_0};
  /* fpexpbf16.vhdl:1086:103  */
  assign n257 = {n256, bh9_w2_0};
  /* fpexpbf16.vhdl:1086:114  */
  assign n258 = {n257, bh9_w1_0};
  /* fpexpbf16.vhdl:1086:125  */
  assign n259 = {n258, bh9_w0_0};
  /* fpexpbf16.vhdl:1089:4  */
  intadder_12_freq500_uid18 bitheapfinaladd_bh9 (
    .clk(clk),
    .x(bitheapfinaladd_bh9_in0),
    .y(bitheapfinaladd_bh9_in1),
    .cin(bitheapfinaladd_bh9_cin),
    .r(bitheapfinaladd_bh9_n261));
  /* fpexpbf16.vhdl:1097:15  */
  assign n264 = outres[11:4]; // extract
endmodule

module intadder_17_freq500_uid38
  (input  clk,
   input  [16:0] x,
   input  [16:0] y,
   input  cin,
   output [16:0] r);
  wire [16:0] rtmp;
  wire [16:0] n209;
  wire [16:0] n210;
  wire [16:0] n211;
  assign r = rtmp; //(module output)
  /* fpexpbf16.vhdl:1554:8  */
  assign rtmp = n211; // (signal)
  /* fpexpbf16.vhdl:1557:14  */
  assign n209 = x + y;
  /* fpexpbf16.vhdl:1557:18  */
  assign n210 = {16'b0, cin};  //  uext
  /* fpexpbf16.vhdl:1557:18  */
  assign n211 = n209 + n210;
endmodule

module exp_8_7_freq500_uid6
  (input  clk,
   input  [15:0] ufixx_i,
   input  xsign,
   output [11:0] expy,
   output [8:0] k);
  wire [15:0] ufixx;
  wire [9:0] xmulin;
  wire [7:0] absk;
  wire [7:0] absk_d1;
  wire [8:0] minusabsk;
  wire [16:0] absklog2;
  wire [8:0] subop1;
  wire [8:0] subop2;
  wire [8:0] y;
  wire xsign_d1;
  wire xsign_d2;
  wire xsign_d3;
  wire [9:0] n174;
  wire [7:0] mulinvlog2_n175;
  wire [8:0] n179;
  wire [8:0] n181;
  wire [8:0] n182;
  wire [8:0] n184;
  wire [16:0] mullog2_n185;
  wire [8:0] n188;
  wire n189;
  wire [8:0] n190;
  wire [8:0] n191;
  wire [8:0] n192;
  wire [8:0] n193;
  wire [8:0] n194;
  wire [8:0] n195;
  wire [8:0] n196;
  localparam n197 = 1'b1;
  wire [8:0] theyadder_n198;
  wire [11:0] expytable_n201;
  reg [7:0] n204;
  reg n205;
  reg n206;
  reg n207;
  assign expy = expytable_n201; //(module output)
  assign k = n182; //(module output)
  /* fpexpbf16.vhdl:1466:8  */
  assign xmulin = n174; // (signal)
  /* fpexpbf16.vhdl:1468:8  */
  assign absk = mulinvlog2_n175; // (signal)
  /* fpexpbf16.vhdl:1468:14  */
  assign absk_d1 = n204; // (signal)
  /* fpexpbf16.vhdl:1470:8  */
  assign minusabsk = n181; // (signal)
  /* fpexpbf16.vhdl:1472:8  */
  assign absklog2 = mullog2_n185; // (signal)
  /* fpexpbf16.vhdl:1474:8  */
  assign subop1 = n190; // (signal)
  /* fpexpbf16.vhdl:1476:8  */
  assign subop2 = n194; // (signal)
  /* fpexpbf16.vhdl:1478:8  */
  assign y = theyadder_n198; // (signal)
  /* fpexpbf16.vhdl:1480:8  */
  assign xsign_d1 = n205; // (signal)
  /* fpexpbf16.vhdl:1480:18  */
  assign xsign_d2 = n206; // (signal)
  /* fpexpbf16.vhdl:1480:28  */
  assign xsign_d3 = n207; // (signal)
  /* fpexpbf16.vhdl:1497:19  */
  assign n174 = ufixx[15:6]; // extract
  /* fpexpbf16.vhdl:1498:4  */
  fixrealkcm_freq500_uid8 mulinvlog2 (
    .clk(clk),
    .x(xmulin),
    .r(mulinvlog2_n175));
  /* fpexpbf16.vhdl:1502:44  */
  assign n179 = {1'b0, absk_d1};
  /* fpexpbf16.vhdl:1502:37  */
  assign n181 = 9'b000000000 - n179;
  /* fpexpbf16.vhdl:1503:19  */
  assign n182 = xsign_d3 ? minusabsk : n184;
  /* fpexpbf16.vhdl:1503:50  */
  assign n184 = {1'b0, absk_d1};
  /* fpexpbf16.vhdl:1504:4  */
  fixrealkcm_freq500_uid20 mullog2 (
    .clk(clk),
    .x(absk),
    .r(mullog2_n185));
  /* fpexpbf16.vhdl:1508:36  */
  assign n188 = ufixx[8:0]; // extract
  /* fpexpbf16.vhdl:1508:63  */
  assign n189 = ~xsign_d1;
  /* fpexpbf16.vhdl:1508:50  */
  assign n190 = n189 ? n188 : n192;
  /* fpexpbf16.vhdl:1508:100  */
  assign n191 = ufixx[8:0]; // extract
  /* fpexpbf16.vhdl:1508:73  */
  assign n192 = ~n191;
  /* fpexpbf16.vhdl:1509:22  */
  assign n193 = absklog2[8:0]; // extract
  /* fpexpbf16.vhdl:1509:35  */
  assign n194 = xsign_d3 ? n193 : n196;
  /* fpexpbf16.vhdl:1509:71  */
  assign n195 = absklog2[8:0]; // extract
  /* fpexpbf16.vhdl:1509:58  */
  assign n196 = ~n195;
  /* fpexpbf16.vhdl:1510:4  */
  intadder_9_freq500_uid33 theyadder (
    .clk(clk),
    .x(subop1),
    .y(subop2),
    .cin(n197),
    .r(theyadder_n198));
  /* fpexpbf16.vhdl:1517:4  */
  fixfunctionbytable_freq500_uid35 expytable (
    .x(y),
    .y(expytable_n201));
  /* fpexpbf16.vhdl:1489:10  */
  always @(posedge clk)
    n204 <= absk;
  /* fpexpbf16.vhdl:1489:10  */
  always @(posedge clk)
    n205 <= xsign;
  /* fpexpbf16.vhdl:1489:10  */
  always @(posedge clk)
    n206 <= xsign_d1;
  /* fpexpbf16.vhdl:1489:10  */
  always @(posedge clk)
    n207 <= xsign_d2;
endmodule

module leftshifter8_by_max_15_freq500_uid4
  (input  clk,
   input  [7:0] x,
   input  [3:0] s,
   output [22:0] r);
  wire [3:0] ps;
  wire [3:0] ps_d1;
  wire [7:0] level0;
  wire [8:0] level1;
  wire [8:0] level1_d1;
  wire [10:0] level2;
  wire [14:0] level3;
  wire [22:0] level4;
  wire [8:0] n139;
  wire n140;
  wire [8:0] n141;
  wire [8:0] n143;
  wire [10:0] n145;
  wire n146;
  wire [10:0] n147;
  wire [10:0] n149;
  wire [14:0] n151;
  wire n152;
  wire [14:0] n153;
  wire [14:0] n155;
  wire [22:0] n157;
  wire n158;
  wire [22:0] n159;
  wire [22:0] n161;
  reg [3:0] n162;
  reg [8:0] n163;
  assign r = level4; //(module output)
  /* fpexpbf16.vhdl:850:12  */
  assign ps_d1 = n162; // (signal)
  /* fpexpbf16.vhdl:854:8  */
  assign level1 = n141; // (signal)
  /* fpexpbf16.vhdl:854:16  */
  assign level1_d1 = n163; // (signal)
  /* fpexpbf16.vhdl:856:8  */
  assign level2 = n147; // (signal)
  /* fpexpbf16.vhdl:858:8  */
  assign level3 = n153; // (signal)
  /* fpexpbf16.vhdl:860:8  */
  assign level4 = n159; // (signal)
  /* fpexpbf16.vhdl:872:20  */
  assign n139 = {level0, 1'b0};
  /* fpexpbf16.vhdl:872:49  */
  assign n140 = ps[0]; // extract
  /* fpexpbf16.vhdl:872:42  */
  assign n141 = n140 ? n139 : n143;
  /* fpexpbf16.vhdl:872:87  */
  assign n143 = {1'b0, level0};
  /* fpexpbf16.vhdl:873:23  */
  assign n145 = {level1_d1, 2'b00};
  /* fpexpbf16.vhdl:873:55  */
  assign n146 = ps_d1[1]; // extract
  /* fpexpbf16.vhdl:873:45  */
  assign n147 = n146 ? n145 : n149;
  /* fpexpbf16.vhdl:873:93  */
  assign n149 = {2'b00, level1_d1};
  /* fpexpbf16.vhdl:874:20  */
  assign n151 = {level2, 4'b0000};
  /* fpexpbf16.vhdl:874:52  */
  assign n152 = ps_d1[2]; // extract
  /* fpexpbf16.vhdl:874:42  */
  assign n153 = n152 ? n151 : n155;
  /* fpexpbf16.vhdl:874:90  */
  assign n155 = {4'b0000, level2};
  /* fpexpbf16.vhdl:875:20  */
  assign n157 = {level3, 8'b00000000};
  /* fpexpbf16.vhdl:875:52  */
  assign n158 = ps_d1[3]; // extract
  /* fpexpbf16.vhdl:875:42  */
  assign n159 = n158 ? n157 : n161;
  /* fpexpbf16.vhdl:875:90  */
  assign n161 = {8'b00000000, level3};
  /* fpexpbf16.vhdl:865:10  */
  always @(posedge clk)
    n162 <= ps;
  /* fpexpbf16.vhdl:865:10  */
  always @(posedge clk)
    n163 <= level1;
endmodule

module top_module
  (input  clk,
   input  [17:0] X,
   output [17:0] R);
  wire [1:0] xexn;
  wire [1:0] xexn_d1;
  wire xsign;
  wire xsign_d1;
  wire [7:0] xexpfield;
  wire [6:0] xfrac;
  wire [9:0] e0;
  wire [9:0] shiftval;
  wire [9:0] shiftval_d1;
  wire resultwillbeone;
  wire resultwillbeone_d1;
  wire [7:0] mxu;
  wire [8:0] maxshift;
  wire [8:0] maxshift_d1;
  wire overflow0;
  wire [3:0] shiftvalin;
  wire [22:0] fixx0;
  wire [15:0] ufixx;
  wire [11:0] expy;
  wire [8:0] k;
  wire neednonorm;
  wire [16:0] preroundbiassig;
  wire roundbit;
  wire [16:0] roundnormaddend;
  wire [16:0] roundedexpsigres;
  wire [16:0] roundedexpsig;
  wire ofl1;
  wire ofl2;
  wire ofl3;
  wire ofl;
  wire ufl1;
  wire ufl2;
  wire ufl3;
  wire ufl;
  wire [1:0] rexn;
  wire [1:0] n10;
  wire n11;
  wire [7:0] n12;
  wire [6:0] n13;
  wire [9:0] n16;
  wire [9:0] n17;
  wire n18;
  wire [7:0] n20;
  wire n22;
  wire n23;
  wire [8:0] n24;
  wire n25;
  wire n26;
  wire [3:0] n28;
  wire [22:0] mantissa_shift_n29;
  wire [15:0] n32;
  wire n33;
  wire [15:0] n34;
  wire [11:0] exp_helper_n36;
  wire [8:0] exp_helper_n37;
  wire n42;
  wire [6:0] n43;
  wire [16:0] n45;
  wire [16:0] n46;
  wire [6:0] n47;
  wire [16:0] n49;
  wire n50;
  wire n51;
  wire n52;
  wire n53;
  wire [9:0] n54;
  wire [15:0] n56;
  wire [16:0] n57;
  localparam n58 = 1'b0;
  wire [16:0] roundedexpsigoperandadder_n59;
  wire n63;
  wire [16:0] n64;
  wire n66;
  wire n67;
  wire n68;
  wire n69;
  wire n70;
  wire n71;
  wire n72;
  wire n73;
  wire n74;
  wire n75;
  wire n76;
  wire n77;
  wire n78;
  wire n79;
  wire n80;
  wire n81;
  wire n82;
  wire n83;
  wire n84;
  wire n85;
  wire n86;
  wire n87;
  wire n88;
  wire n89;
  wire n90;
  wire n91;
  wire n92;
  wire n93;
  wire n94;
  wire n95;
  wire n96;
  wire n97;
  wire n98;
  wire n99;
  wire n100;
  wire n101;
  wire n102;
  wire n103;
  wire n104;
  wire n105;
  wire n106;
  wire n107;
  wire n108;
  wire n109;
  wire n110;
  wire n111;
  wire n112;
  wire n115;
  wire [1:0] n116;
  wire [1:0] n118;
  wire [1:0] n120;
  wire [2:0] n123;
  wire [14:0] n124;
  wire [17:0] n125;
  reg [1:0] n126;
  reg n127;
  reg [9:0] n128;
  reg n129;
  reg [8:0] n130;
  assign R = n125; //(module output)
  /* fpexpbf16.vhdl:1615:8  */
  assign xexn = n10; // (signal)
  /* fpexpbf16.vhdl:1615:14  */
  assign xexn_d1 = n126; // (signal)
  /* fpexpbf16.vhdl:1617:8  */
  assign xsign = n11; // (signal)
  /* fpexpbf16.vhdl:1617:15  */
  assign xsign_d1 = n127; // (signal)
  /* fpexpbf16.vhdl:1619:8  */
  assign xexpfield = n12; // (signal)
  /* fpexpbf16.vhdl:1621:8  */
  assign xfrac = n13; // (signal)
  /* fpexpbf16.vhdl:1623:8  */
  assign e0 = 10'b0001110110; // (signal)
  /* fpexpbf16.vhdl:1625:8  */
  assign shiftval = n17; // (signal)
  /* fpexpbf16.vhdl:1625:18  */
  assign shiftval_d1 = n128; // (signal)
  /* fpexpbf16.vhdl:1627:8  */
  assign resultwillbeone = n18; // (signal)
  /* fpexpbf16.vhdl:1627:25  */
  assign resultwillbeone_d1 = n129; // (signal)
  /* fpexpbf16.vhdl:1629:8  */
  assign mxu = n20; // (signal)
  /* fpexpbf16.vhdl:1631:8  */
  assign maxshift = 9'b000001111; // (signal)
  /* fpexpbf16.vhdl:1631:18  */
  assign maxshift_d1 = n130; // (signal)
  /* fpexpbf16.vhdl:1633:8  */
  assign overflow0 = n26; // (signal)
  /* fpexpbf16.vhdl:1635:8  */
  assign shiftvalin = n28; // (signal)
  /* fpexpbf16.vhdl:1637:8  */
  assign fixx0 = mantissa_shift_n29; // (signal)
  /* fpexpbf16.vhdl:1639:8  */
  assign ufixx = n34; // (signal)
  /* fpexpbf16.vhdl:1641:8  */
  assign expy = exp_helper_n36; // (signal)
  /* fpexpbf16.vhdl:1643:8  */
  assign k = exp_helper_n37; // (signal)
  /* fpexpbf16.vhdl:1645:8  */
  assign neednonorm = n42; // (signal)
  /* fpexpbf16.vhdl:1647:8  */
  assign preroundbiassig = n46; // (signal)
  /* fpexpbf16.vhdl:1649:8  */
  assign roundbit = n51; // (signal)
  /* fpexpbf16.vhdl:1651:8  */
  assign roundnormaddend = n57; // (signal)
  /* fpexpbf16.vhdl:1653:8  */
  assign roundedexpsigres = roundedexpsigoperandadder_n59; // (signal)
  /* fpexpbf16.vhdl:1655:8  */
  assign roundedexpsig = n64; // (signal)
  /* fpexpbf16.vhdl:1657:8  */
  assign ofl1 = n72; // (signal)
  /* fpexpbf16.vhdl:1659:8  */
  assign ofl2 = n83; // (signal)
  /* fpexpbf16.vhdl:1661:8  */
  assign ofl3 = n89; // (signal)
  /* fpexpbf16.vhdl:1663:8  */
  assign ofl = n91; // (signal)
  /* fpexpbf16.vhdl:1665:8  */
  assign ufl1 = n99; // (signal)
  /* fpexpbf16.vhdl:1667:8  */
  assign ufl2 = n104; // (signal)
  /* fpexpbf16.vhdl:1669:8  */
  assign ufl3 = n110; // (signal)
  /* fpexpbf16.vhdl:1671:8  */
  assign ufl = n112; // (signal)
  /* fpexpbf16.vhdl:1673:8  */
  assign rexn = n116; // (signal)
  /* fpexpbf16.vhdl:1690:13  */
  assign n10 = X[17:16]; // extract
  /* fpexpbf16.vhdl:1691:14  */
  assign n11 = X[15]; // extract
  /* fpexpbf16.vhdl:1692:18  */
  assign n12 = X[14:7]; // extract
  /* fpexpbf16.vhdl:1693:23  */
  assign n13 = X[6:0]; // extract
  /* fpexpbf16.vhdl:1695:22  */
  assign n16 = {2'b00, xexpfield};
  /* fpexpbf16.vhdl:1695:35  */
  assign n17 = n16 - e0;
  /* fpexpbf16.vhdl:1697:31  */
  assign n18 = shiftval[9]; // extract
  /* fpexpbf16.vhdl:1699:15  */
  assign n20 = {1'b1, xfrac};
  /* fpexpbf16.vhdl:1702:32  */
  assign n22 = shiftval_d1[9]; // extract
  /* fpexpbf16.vhdl:1702:17  */
  assign n23 = ~n22;
  /* fpexpbf16.vhdl:1702:55  */
  assign n24 = shiftval_d1[8:0]; // extract
  /* fpexpbf16.vhdl:1702:69  */
  assign n25 = $unsigned(n24) > $unsigned(maxshift_d1);
  /* fpexpbf16.vhdl:1702:39  */
  assign n26 = n25 ? n23 : 1'b0;
  /* fpexpbf16.vhdl:1703:26  */
  assign n28 = shiftval[3:0]; // extract
  /* fpexpbf16.vhdl:1704:4  */
  leftshifter8_by_max_15_freq500_uid4 mantissa_shift (
    .clk(clk),
    .x(mxu),
    .s(shiftvalin),
    .r(mantissa_shift_n29));
  /* fpexpbf16.vhdl:1709:28  */
  assign n32 = fixx0[22:7]; // extract
  /* fpexpbf16.vhdl:1709:66  */
  assign n33 = ~resultwillbeone_d1;
  /* fpexpbf16.vhdl:1709:43  */
  assign n34 = n33 ? n32 : 16'b0000000000000000;
  /* fpexpbf16.vhdl:1710:4  */
  exp_8_7_freq500_uid6 exp_helper (
    .clk(clk),
    .ufixx_i(ufixx),
    .xsign(xsign),
    .expy(exp_helper_n36),
    .k(exp_helper_n37));
  /* fpexpbf16.vhdl:1716:22  */
  assign n42 = expy[11]; // extract
  /* fpexpbf16.vhdl:1718:63  */
  assign n43 = expy[10:4]; // extract
  /* fpexpbf16.vhdl:1718:57  */
  assign n45 = {10'b0001111111, n43};
  /* fpexpbf16.vhdl:1718:77  */
  assign n46 = neednonorm ? n45 : n49;
  /* fpexpbf16.vhdl:1719:52  */
  assign n47 = expy[9:3]; // extract
  /* fpexpbf16.vhdl:1719:46  */
  assign n49 = {10'b0001111110, n47};
  /* fpexpbf16.vhdl:1720:20  */
  assign n50 = expy[3]; // extract
  /* fpexpbf16.vhdl:1720:25  */
  assign n51 = neednonorm ? n50 : n52;
  /* fpexpbf16.vhdl:1720:59  */
  assign n52 = expy[2]; // extract
  /* fpexpbf16.vhdl:1721:24  */
  assign n53 = k[8]; // extract
  /* fpexpbf16.vhdl:1721:28  */
  assign n54 = {n53, k};
  /* fpexpbf16.vhdl:1721:32  */
  assign n56 = {n54, 6'b000000};
  /* fpexpbf16.vhdl:1721:54  */
  assign n57 = {n56, roundbit};
  /* fpexpbf16.vhdl:1722:4  */
  intadder_17_freq500_uid38 roundedexpsigoperandadder (
    .clk(clk),
    .x(preroundbiassig),
    .y(roundnormaddend),
    .cin(n58),
    .r(roundedexpsigoperandadder_n59));
  /* fpexpbf16.vhdl:1728:47  */
  assign n63 = xexn == 2'b01;
  /* fpexpbf16.vhdl:1728:38  */
  assign n64 = n63 ? roundedexpsigres : 17'b00011111110000000;
  /* fpexpbf16.vhdl:1729:12  */
  assign n66 = ~xsign_d1;
  /* fpexpbf16.vhdl:1729:25  */
  assign n67 = n66 & overflow0;
  /* fpexpbf16.vhdl:1729:55  */
  assign n68 = xexn_d1[1]; // extract
  /* fpexpbf16.vhdl:1729:44  */
  assign n69 = ~n68;
  /* fpexpbf16.vhdl:1729:70  */
  assign n70 = xexn_d1[0]; // extract
  /* fpexpbf16.vhdl:1729:59  */
  assign n71 = n69 & n70;
  /* fpexpbf16.vhdl:1729:39  */
  assign n72 = n67 & n71;
  /* fpexpbf16.vhdl:1730:12  */
  assign n73 = ~xsign;
  /* fpexpbf16.vhdl:1730:40  */
  assign n74 = roundedexpsig[15]; // extract
  /* fpexpbf16.vhdl:1730:69  */
  assign n75 = roundedexpsig[16]; // extract
  /* fpexpbf16.vhdl:1730:52  */
  assign n76 = ~n75;
  /* fpexpbf16.vhdl:1730:48  */
  assign n77 = n74 & n76;
  /* fpexpbf16.vhdl:1730:22  */
  assign n78 = n73 & n77;
  /* fpexpbf16.vhdl:1730:93  */
  assign n79 = xexn[1]; // extract
  /* fpexpbf16.vhdl:1730:85  */
  assign n80 = ~n79;
  /* fpexpbf16.vhdl:1730:105  */
  assign n81 = xexn[0]; // extract
  /* fpexpbf16.vhdl:1730:97  */
  assign n82 = n80 & n81;
  /* fpexpbf16.vhdl:1730:80  */
  assign n83 = n78 & n82;
  /* fpexpbf16.vhdl:1731:12  */
  assign n84 = ~xsign;
  /* fpexpbf16.vhdl:1731:30  */
  assign n85 = xexn[1]; // extract
  /* fpexpbf16.vhdl:1731:22  */
  assign n86 = n84 & n85;
  /* fpexpbf16.vhdl:1731:46  */
  assign n87 = xexn[0]; // extract
  /* fpexpbf16.vhdl:1731:38  */
  assign n88 = ~n87;
  /* fpexpbf16.vhdl:1731:34  */
  assign n89 = n86 & n88;
  /* fpexpbf16.vhdl:1732:16  */
  assign n90 = ofl1 | ofl2;
  /* fpexpbf16.vhdl:1732:24  */
  assign n91 = n90 | ofl3;
  /* fpexpbf16.vhdl:1733:26  */
  assign n92 = roundedexpsig[15]; // extract
  /* fpexpbf16.vhdl:1733:51  */
  assign n93 = roundedexpsig[16]; // extract
  /* fpexpbf16.vhdl:1733:34  */
  assign n94 = n92 & n93;
  /* fpexpbf16.vhdl:1733:76  */
  assign n95 = xexn[1]; // extract
  /* fpexpbf16.vhdl:1733:68  */
  assign n96 = ~n95;
  /* fpexpbf16.vhdl:1733:88  */
  assign n97 = xexn[0]; // extract
  /* fpexpbf16.vhdl:1733:80  */
  assign n98 = n96 & n97;
  /* fpexpbf16.vhdl:1733:63  */
  assign n99 = n94 & n98;
  /* fpexpbf16.vhdl:1734:26  */
  assign n100 = xexn[1]; // extract
  /* fpexpbf16.vhdl:1734:18  */
  assign n101 = xsign & n100;
  /* fpexpbf16.vhdl:1734:42  */
  assign n102 = xexn[0]; // extract
  /* fpexpbf16.vhdl:1734:34  */
  assign n103 = ~n102;
  /* fpexpbf16.vhdl:1734:30  */
  assign n104 = n101 & n103;
  /* fpexpbf16.vhdl:1735:21  */
  assign n105 = xsign_d1 & overflow0;
  /* fpexpbf16.vhdl:1735:52  */
  assign n106 = xexn_d1[1]; // extract
  /* fpexpbf16.vhdl:1735:41  */
  assign n107 = ~n106;
  /* fpexpbf16.vhdl:1735:67  */
  assign n108 = xexn_d1[0]; // extract
  /* fpexpbf16.vhdl:1735:56  */
  assign n109 = n107 & n108;
  /* fpexpbf16.vhdl:1735:36  */
  assign n110 = n105 & n109;
  /* fpexpbf16.vhdl:1736:16  */
  assign n111 = ufl1 | ufl2;
  /* fpexpbf16.vhdl:1736:24  */
  assign n112 = n111 | ufl3;
  /* fpexpbf16.vhdl:1737:27  */
  assign n115 = xexn == 2'b11;
  /* fpexpbf16.vhdl:1737:17  */
  assign n116 = n115 ? 2'b11 : n118;
  /* fpexpbf16.vhdl:1738:7  */
  assign n118 = ofl ? 2'b10 : n120;
  /* fpexpbf16.vhdl:1739:7  */
  assign n120 = ufl ? 2'b00 : 2'b01;
  /* fpexpbf16.vhdl:1741:14  */
  assign n123 = {rexn, 1'b0};
  /* fpexpbf16.vhdl:1741:35  */
  assign n124 = roundedexpsig[14:0]; // extract
  /* fpexpbf16.vhdl:1741:20  */
  assign n125 = {n123, n124};
  /* fpexpbf16.vhdl:1682:10  */
  always @(posedge clk)
    n126 <= xexn;
  /* fpexpbf16.vhdl:1682:10  */
  always @(posedge clk)
    n127 <= xsign;
  /* fpexpbf16.vhdl:1682:10  */
  always @(posedge clk)
    n128 <= shiftval;
  /* fpexpbf16.vhdl:1682:10  */
  always @(posedge clk)
    n129 <= resultwillbeone;
  /* fpexpbf16.vhdl:1682:10  */
  always @(posedge clk)
    n130 <= maxshift;
endmodule

