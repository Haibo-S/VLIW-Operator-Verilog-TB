--------------------------------------------------------------------------------
--                          InvA0Table_Freq500_uid15
-- VHDL generated for DummyFPGA @ 500MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 2
-- Target frequency (MHz): 500
-- Input signals: X
-- Output signals: Y
--  approx. input signal timings: X: (c0, 0.000000ns)
--  approx. output signal timings: Y: (c0, 0.550000ns)

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity InvA0Table_Freq500_uid15 is
    port (X : in  std_logic_vector(6 downto 0);
          Y : out  std_logic_vector(7 downto 0)   );
end entity;

architecture arch of InvA0Table_Freq500_uid15 is
signal Y0 :  std_logic_vector(7 downto 0);
   -- timing of Y0: (c0, 0.550000ns)
signal Y1 :  std_logic_vector(7 downto 0);
   -- timing of Y1: (c0, 0.550000ns)
begin
   with X  select  Y0 <= 
      "10000000" when "0000000",
      "10000000" when "0000001",
      "01111111" when "0000010",
      "01111110" when "0000011",
      "01111101" when "0000100",
      "01111100" when "0000101",
      "01111011" when "0000110",
      "01111010" when "0000111",
      "01111001" when "0001000",
      "01111000" when "0001001",
      "01110111" when "0001010",
      "01110110" when "0001011",
      "01110110" when "0001100",
      "01110101" when "0001101",
      "01110100" when "0001110",
      "01110011" when "0001111",
      "01110010" when "0010000",
      "01110001" when "0010001",
      "01110001" when "0010010",
      "01110000" when "0010011",
      "01101111" when "0010100",
      "01101110" when "0010101",
      "01101110" when "0010110",
      "01101101" when "0010111",
      "01101100" when "0011000",
      "01101100" when "0011001",
      "01101011" when "0011010",
      "01101010" when "0011011",
      "01101010" when "0011100",
      "01101001" when "0011101",
      "01101000" when "0011110",
      "01101000" when "0011111",
      "01100111" when "0100000",
      "01100110" when "0100001",
      "01100110" when "0100010",
      "01100101" when "0100011",
      "01100100" when "0100100",
      "01100100" when "0100101",
      "01100011" when "0100110",
      "01100011" when "0100111",
      "01100010" when "0101000",
      "01100001" when "0101001",
      "01100001" when "0101010",
      "01100000" when "0101011",
      "01100000" when "0101100",
      "01011111" when "0101101",
      "01011111" when "0101110",
      "01011110" when "0101111",
      "01011110" when "0110000",
      "01011101" when "0110001",
      "01011101" when "0110010",
      "01011100" when "0110011",
      "01011100" when "0110100",
      "01011011" when "0110101",
      "01011011" when "0110110",
      "01011010" when "0110111",
      "01011010" when "0111000",
      "01011001" when "0111001",
      "01011001" when "0111010",
      "01011000" when "0111011",
      "01011000" when "0111100",
      "01010111" when "0111101",
      "01010111" when "0111110",
      "01010110" when "0111111",
      "10101011" when "1000000",
      "10101010" when "1000001",
      "10101001" when "1000010",
      "10101001" when "1000011",
      "10101000" when "1000100",
      "10100111" when "1000101",
      "10100110" when "1000110",
      "10100101" when "1000111",
      "10100100" when "1001000",
      "10100100" when "1001001",
      "10100011" when "1001010",
      "10100010" when "1001011",
      "10100001" when "1001100",
      "10100000" when "1001101",
      "10100000" when "1001110",
      "10011111" when "1001111",
      "10011110" when "1010000",
      "10011101" when "1010001",
      "10011101" when "1010010",
      "10011100" when "1010011",
      "10011011" when "1010100",
      "10011010" when "1010101",
      "10011010" when "1010110",
      "10011001" when "1010111",
      "10011000" when "1011000",
      "10011000" when "1011001",
      "10010111" when "1011010",
      "10010110" when "1011011",
      "10010101" when "1011100",
      "10010101" when "1011101",
      "10010100" when "1011110",
      "10010011" when "1011111",
      "10010011" when "1100000",
      "10010010" when "1100001",
      "10010001" when "1100010",
      "10010001" when "1100011",
      "10010000" when "1100100",
      "10010000" when "1100101",
      "10001111" when "1100110",
      "10001110" when "1100111",
      "10001110" when "1101000",
      "10001101" when "1101001",
      "10001101" when "1101010",
      "10001100" when "1101011",
      "10001011" when "1101100",
      "10001011" when "1101101",
      "10001010" when "1101110",
      "10001010" when "1101111",
      "10001001" when "1110000",
      "10001000" when "1110001",
      "10001000" when "1110010",
      "10000111" when "1110011",
      "10000111" when "1110100",
      "10000110" when "1110101",
      "10000110" when "1110110",
      "10000101" when "1110111",
      "10000101" when "1111000",
      "10000100" when "1111001",
      "10000100" when "1111010",
      "10000011" when "1111011",
      "10000011" when "1111100",
      "10000010" when "1111101",
      "10000010" when "1111110",
      "10000001" when "1111111",
      "--------" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          LogTable0_Freq500_uid27
-- VHDL generated for DummyFPGA @ 500MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 2
-- Target frequency (MHz): 500
-- Input signals: X
-- Output signals: Y
--  approx. input signal timings: X: (c0, 0.000000ns)
--  approx. output signal timings: Y: (c0, 0.550000ns)

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity LogTable0_Freq500_uid27 is
    port (X : in  std_logic_vector(6 downto 0);
          Y : out  std_logic_vector(29 downto 0)   );
end entity;

architecture arch of LogTable0_Freq500_uid27 is
signal Y0 :  std_logic_vector(29 downto 0);
   -- timing of Y0: (c0, 0.550000ns)
signal Y1 :  std_logic_vector(29 downto 0);
   -- timing of Y1: (c0, 0.550000ns)
begin
   with X  select  Y0 <= 
      "111111111100000000000000000000" when "0000000",
      "111111111100000000000000000000" when "0000001",
      "000000011100001000000010101100" when "0000010",
      "000000111100100000010101100110" when "0000011",
      "000001011101001001001001010011" when "0000100",
      "000001111110000010101110110001" when "0000101",
      "000010011111001101010111011010" when "0000110",
      "000011000000101001010101000011" when "0000111",
      "000011100010010110111001111010" when "0001000",
      "000100000100010110011000101101" when "0001001",
      "000100100110101000000100101001" when "0001010",
      "000101001001001100010001010111" when "0001011",
      "000101001001001100010001010111" when "0001100",
      "000101101100000011010011000011" when "0001101",
      "000110001111001101011110010111" when "0001110",
      "000110110010101011001000100011" when "0001111",
      "000111010110011100100111011001" when "0010000",
      "000111111010100010010001001110" when "0010001",
      "000111111010100010010001001110" when "0010010",
      "001000011110111100011101000001" when "0010011",
      "001001000011101011100010010101" when "0010100",
      "001001101000101111111001011000" when "0010101",
      "001001101000101111111001011000" when "0010110",
      "001010001110001001111011000010" when "0010111",
      "001010110011111010000000110110" when "0011000",
      "001010110011111010000000110110" when "0011001",
      "001011011010000000100101000110" when "0011010",
      "001100000000011110000010110011" when "0011011",
      "001100000000011110000010110011" when "0011100",
      "001100100111010010110101101110" when "0011101",
      "001101001110011111011010011110" when "0011110",
      "001101001110011111011010011110" when "0011111",
      "001101110110000100001110011100" when "0100000",
      "001110011110000001101111111001" when "0100001",
      "001110011110000001101111111001" when "0100010",
      "001111000110011000011110000000" when "0100011",
      "001111101111001000111000110110" when "0100100",
      "001111101111001000111000110110" when "0100101",
      "010000011000010011100001100000" when "0100110",
      "010000011000010011100001100000" when "0100111",
      "010001000001111000111010000010" when "0101000",
      "010001101011111001100101100100" when "0101001",
      "010001101011111001100101100100" when "0101010",
      "010010010110010110001000010001" when "0101011",
      "010010010110010110001000010001" when "0101100",
      "010011000001001111000111100010" when "0101101",
      "010011000001001111000111100010" when "0101110",
      "010011101100100101001001110111" when "0101111",
      "010011101100100101001001110111" when "0110000",
      "010100011000011000110111000010" when "0110001",
      "010100011000011000110111000010" when "0110010",
      "010101000100101010111000000111" when "0110011",
      "010101000100101010111000000111" when "0110100",
      "010101110001011011110111100000" when "0110101",
      "010101110001011011110111100000" when "0110110",
      "010110011110101100100000111110" when "0110111",
      "010110011110101100100000111110" when "0111000",
      "010111001100011101100001110111" when "0111001",
      "010111001100011101100001110111" when "0111010",
      "010111111010101111101000111100" when "0111011",
      "010111111010101111101000111100" when "0111100",
      "011000101001100011100110101000" when "0111101",
      "011000101001100011100110101000" when "0111110",
      "011001011000111010001101000011" when "0111111",
      "101101011001101010010111101100" when "1000000",
      "101101110001101011111000000100" when "1000001",
      "101110001001110110011100111110" when "1000010",
      "101110001001110110011100111110" when "1000011",
      "101110100010001010001101010100" when "1000100",
      "101110111010100111010000000110" when "1000101",
      "101111010011001101101100011110" when "1000110",
      "101111101011111101101001101100" when "1000111",
      "110000000100110111001111001001" when "1001000",
      "110000000100110111001111001001" when "1001001",
      "110000011101111010100100011010" when "1001010",
      "110000110111000111110001001001" when "1001011",
      "110001010000011110111101001010" when "1001100",
      "110001101010000000010000011100" when "1001101",
      "110001101010000000010000011100" when "1001110",
      "110010000011101011110011000110" when "1001111",
      "110010011101100001101101011001" when "1010000",
      "110010110111100010000111110000" when "1010001",
      "110010110111100010000111110000" when "1010010",
      "110011010001101101001010110010" when "1010011",
      "110011101100000010111111001110" when "1010100",
      "110100000110100011101101111111" when "1010101",
      "110100000110100011101101111111" when "1010110",
      "110100100001001111100000001100" when "1010111",
      "110100111100000110011111001000" when "1011000",
      "110100111100000110011111001000" when "1011001",
      "110101010111001000110100001110" when "1011010",
      "110101110010010110101001001010" when "1011011",
      "110110001101110000000111110000" when "1011100",
      "110110001101110000000111110000" when "1011101",
      "110110101001010101011010000100" when "1011110",
      "110111000101000110101010010110" when "1011111",
      "110111000101000110101010010110" when "1100000",
      "110111100001000100000011000010" when "1100001",
      "110111111101001101101110110100" when "1100010",
      "110111111101001101101110110100" when "1100011",
      "111000011001100011111000100100" when "1100100",
      "111000011001100011111000100100" when "1100101",
      "111000110110000110101011011100" when "1100110",
      "111001010010110110010010110001" when "1100111",
      "111001010010110110010010110001" when "1101000",
      "111001101111110010111010001010" when "1101001",
      "111001101111110010111010001010" when "1101010",
      "111010001100111100101101011101" when "1101011",
      "111010101010010011111000110000" when "1101100",
      "111010101010010011111000110000" when "1101101",
      "111011000111111000101000011010" when "1101110",
      "111011000111111000101000011010" when "1101111",
      "111011100101101011001001000100" when "1110000",
      "111100000011101011100111101000" when "1110001",
      "111100000011101011100111101000" when "1110010",
      "111100100001111010010001010010" when "1110011",
      "111100100001111010010001010010" when "1110100",
      "111101000000010111010011100001" when "1110101",
      "111101000000010111010011100001" when "1110110",
      "111101011111000010111100001001" when "1110111",
      "111101011111000010111100001001" when "1111000",
      "111101111101111101011001001111" when "1111001",
      "111101111101111101011001001111" when "1111010",
      "111110011101000110111001010000" when "1111011",
      "111110011101000110111001010000" when "1111100",
      "111110111100011111101010111010" when "1111101",
      "111110111100011111101010111010" when "1111110",
      "111111011100000111111101010110" when "1111111",
      "------------------------------" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          LogTable1_Freq500_uid30
-- VHDL generated for DummyFPGA @ 500MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 2
-- Target frequency (MHz): 500
-- Input signals: X
-- Output signals: Y
--  approx. input signal timings: X: (c0, 0.000000ns)
--  approx. output signal timings: Y: (c0, 0.550000ns)

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity LogTable1_Freq500_uid30 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(24 downto 0)   );
end entity;

architecture arch of LogTable1_Freq500_uid30 is
signal Y0 :  std_logic_vector(24 downto 0);
   -- timing of Y0: (c0, 0.550000ns)
signal Y1 :  std_logic_vector(24 downto 0);
   -- timing of Y1: (c0, 0.550000ns)
begin
   with X  select  Y0 <= 
      "0000010000000000010000000" when "00000",
      "0000110000000000010000000" when "00001",
      "0001010000000010010000001" when "00010",
      "0001110000000110010000101" when "00011",
      "0010010000001100010001110" when "00100",
      "0010110000010100010011110" when "00101",
      "0011010000011110010111000" when "00110",
      "0011110000101010011011100" when "00111",
      "0100010000111000100001110" when "01000",
      "0100110001001000101001110" when "01001",
      "0101010001011010110100000" when "01010",
      "0101110001101111000000101" when "01011",
      "0110010010000101010000000" when "01100",
      "0110110010011101100010001" when "01101",
      "0111010010110111110111100" when "01110",
      "0111110011010100010000011" when "01111",
      "1000000011100011001110010" when "10000",
      "1000100100000010101100110" when "10001",
      "1001000100100100001111010" when "10010",
      "1001100101000111110110010" when "10011",
      "1010000101101101100001111" when "10100",
      "1010100110010101010010010" when "10101",
      "1011000110111111000111111" when "10110",
      "1011100111101011000011000" when "10111",
      "1100001000011001000011101" when "11000",
      "1100101001001001001010011" when "11001",
      "1101001001111011010111010" when "11010",
      "1101101010101111101010101" when "11011",
      "1110001011100110000100110" when "11100",
      "1110101100011110100101111" when "11101",
      "1111001101011001001110010" when "11110",
      "1111101110010101111110011" when "11111",
      "-------------------------" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                 FixRealKCM_Freq500_uid39_T0_Freq500_uid42
-- VHDL generated for DummyFPGA @ 500MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 2
-- Target frequency (MHz): 500
-- Input signals: X
-- Output signals: Y
--  approx. input signal timings: X: (c0, 0.000000ns)
--  approx. output signal timings: Y: (c0, 0.550000ns)

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity FixRealKCM_Freq500_uid39_T0_Freq500_uid42 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(28 downto 0)   );
end entity;

architecture arch of FixRealKCM_Freq500_uid39_T0_Freq500_uid42 is
signal Y0 :  std_logic_vector(28 downto 0);
   -- timing of Y0: (c0, 0.550000ns)
signal Y1 :  std_logic_vector(28 downto 0);
   -- timing of Y1: (c0, 0.550000ns)
begin
   with X  select  Y0 <= 
      "00000000000000000000000000000" when "00000",
      "00000101100010111001000011000" when "00001",
      "00001011000101110010000110000" when "00010",
      "00010000101000101011001001000" when "00011",
      "00010110001011100100001100000" when "00100",
      "00011011101110011101001111000" when "00101",
      "00100001010001010110010010000" when "00110",
      "00100110110100001111010101000" when "00111",
      "00101100010111001000011000000" when "01000",
      "00110001111010000001011011000" when "01001",
      "00110111011100111010011110000" when "01010",
      "00111100111111110011100001000" when "01011",
      "01000010100010101100100100000" when "01100",
      "01001000000101100101100111000" when "01101",
      "01001101101000011110101010000" when "01110",
      "01010011001011010111101101000" when "01111",
      "01011000101110010000101111111" when "10000",
      "01011110010001001001110010111" when "10001",
      "01100011110100000010110101111" when "10010",
      "01101001010110111011111000111" when "10011",
      "01101110111001110100111011111" when "10100",
      "01110100011100101101111110111" when "10101",
      "01111001111111100111000001111" when "10110",
      "01111111100010100000000100111" when "10111",
      "10000101000101011001000111111" when "11000",
      "10001010101000010010001010111" when "11001",
      "10010000001011001011001101111" when "11010",
      "10010101101110000100010000111" when "11011",
      "10011011010000111101010011111" when "11100",
      "10100000110011110110010110111" when "11101",
      "10100110010110101111011001111" when "11110",
      "10101011111001101000011100111" when "11111",
      "-----------------------------" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                 FixRealKCM_Freq500_uid39_T1_Freq500_uid45
-- VHDL generated for DummyFPGA @ 500MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 2
-- Target frequency (MHz): 500
-- Input signals: X
-- Output signals: Y
--  approx. input signal timings: X: (c0, 0.000000ns)
--  approx. output signal timings: Y: (c0, 0.550000ns)

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity FixRealKCM_Freq500_uid39_T1_Freq500_uid45 is
    port (X : in  std_logic_vector(2 downto 0);
          Y : out  std_logic_vector(23 downto 0)   );
end entity;

architecture arch of FixRealKCM_Freq500_uid39_T1_Freq500_uid45 is
signal Y0 :  std_logic_vector(23 downto 0);
   -- timing of Y0: (c0, 0.550000ns)
signal Y1 :  std_logic_vector(23 downto 0);
   -- timing of Y1: (c0, 0.550000ns)
begin
   with X  select  Y0 <= 
      "000000000000000000000000" when "000",
      "000101100010111001000011" when "001",
      "001011000101110010000110" when "010",
      "010000101000101011001001" when "011",
      "010110001011100100001100" when "100",
      "011011101110011101001111" when "101",
      "100001010001010110010010" when "110",
      "100110110100001111010101" when "111",
      "------------------------" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                 FixRealKCM_Freq500_uid77_T0_Freq500_uid80
-- VHDL generated for DummyFPGA @ 500MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 2
-- Target frequency (MHz): 500
-- Input signals: X
-- Output signals: Y
--  approx. input signal timings: X: (c0, 0.000000ns)
--  approx. output signal timings: Y: (c0, 0.550000ns)

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity FixRealKCM_Freq500_uid77_T0_Freq500_uid80 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(11 downto 0)   );
end entity;

architecture arch of FixRealKCM_Freq500_uid77_T0_Freq500_uid80 is
signal Y0 :  std_logic_vector(11 downto 0);
   -- timing of Y0: (c0, 0.550000ns)
signal Y1 :  std_logic_vector(11 downto 0);
   -- timing of Y1: (c0, 0.550000ns)
begin
   with X  select  Y0 <= 
      "000000001000" when "00000",
      "000001100100" when "00001",
      "000011000001" when "00010",
      "000100011101" when "00011",
      "000101111001" when "00100",
      "000111010110" when "00101",
      "001000110010" when "00110",
      "001010001110" when "00111",
      "001011101011" when "01000",
      "001101000111" when "01001",
      "001110100011" when "01010",
      "010000000000" when "01011",
      "010001011100" when "01100",
      "010010111000" when "01101",
      "010100010101" when "01110",
      "010101110001" when "01111",
      "010111001101" when "10000",
      "011000101010" when "10001",
      "011010000110" when "10010",
      "011011100010" when "10011",
      "011100111111" when "10100",
      "011110011011" when "10101",
      "011111110111" when "10110",
      "100001010100" when "10111",
      "100010110000" when "11000",
      "100100001100" when "11001",
      "100101101001" when "11010",
      "100111000101" when "11011",
      "101000100001" when "11100",
      "101001111110" when "11101",
      "101011011010" when "11110",
      "101100110110" when "11111",
      "------------" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                 FixRealKCM_Freq500_uid77_T1_Freq500_uid83
-- VHDL generated for DummyFPGA @ 500MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 2
-- Target frequency (MHz): 500
-- Input signals: X
-- Output signals: Y
--  approx. input signal timings: X: (c0, 0.000000ns)
--  approx. output signal timings: Y: (c0, 0.550000ns)

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity FixRealKCM_Freq500_uid77_T1_Freq500_uid83 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(6 downto 0)   );
end entity;

architecture arch of FixRealKCM_Freq500_uid77_T1_Freq500_uid83 is
signal Y0 :  std_logic_vector(6 downto 0);
   -- timing of Y0: (c0, 0.550000ns)
signal Y1 :  std_logic_vector(6 downto 0);
   -- timing of Y1: (c0, 0.550000ns)
begin
   with X  select  Y0 <= 
      "0000000" when "00000",
      "0000011" when "00001",
      "0000110" when "00010",
      "0001001" when "00011",
      "0001100" when "00100",
      "0001110" when "00101",
      "0010001" when "00110",
      "0010100" when "00111",
      "0010111" when "01000",
      "0011010" when "01001",
      "0011101" when "01010",
      "0100000" when "01011",
      "0100011" when "01100",
      "0100110" when "01101",
      "0101000" when "01110",
      "0101011" when "01111",
      "0101110" when "10000",
      "0110001" when "10001",
      "0110100" when "10010",
      "0110111" when "10011",
      "0111010" when "10100",
      "0111101" when "10101",
      "0111111" when "10110",
      "1000010" when "10111",
      "1000101" when "11000",
      "1001000" when "11001",
      "1001011" when "11010",
      "1001110" when "11011",
      "1010001" when "11100",
      "1010100" when "11101",
      "1010111" when "11110",
      "1011001" when "11111",
      "-------" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                 FixRealKCM_Freq500_uid89_T0_Freq500_uid92
-- VHDL generated for DummyFPGA @ 500MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 2
-- Target frequency (MHz): 500
-- Input signals: X
-- Output signals: Y
--  approx. input signal timings: X: (c0, 0.000000ns)
--  approx. output signal timings: Y: (c0, 0.550000ns)

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity FixRealKCM_Freq500_uid89_T0_Freq500_uid92 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(17 downto 0)   );
end entity;

architecture arch of FixRealKCM_Freq500_uid89_T0_Freq500_uid92 is
signal Y0 :  std_logic_vector(17 downto 0);
   -- timing of Y0: (c0, 0.550000ns)
signal Y1 :  std_logic_vector(17 downto 0);
   -- timing of Y1: (c0, 0.550000ns)
begin
   with X  select  Y0 <= 
      "000000000000000000" when "00000",
      "000001011000101110" when "00001",
      "000010110001011101" when "00010",
      "000100001010001011" when "00011",
      "000101100010111001" when "00100",
      "000110111011100111" when "00101",
      "001000010100010110" when "00110",
      "001001101101000100" when "00111",
      "001011000101110010" when "01000",
      "001100011110100000" when "01001",
      "001101110111001111" when "01010",
      "001111001111111101" when "01011",
      "010000101000101011" when "01100",
      "010010000001011001" when "01101",
      "010011011010001000" when "01110",
      "010100110010110110" when "01111",
      "010110001011100100" when "10000",
      "010111100100010010" when "10001",
      "011000111101000001" when "10010",
      "011010010101101111" when "10011",
      "011011101110011101" when "10100",
      "011101000111001011" when "10101",
      "011110011111111010" when "10110",
      "011111111000101000" when "10111",
      "100001010001010110" when "11000",
      "100010101010000101" when "11001",
      "100100000010110011" when "11010",
      "100101011011100001" when "11011",
      "100110110100001111" when "11100",
      "101000001100111110" when "11101",
      "101001100101101100" when "11110",
      "101010111110011010" when "11111",
      "------------------" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                 FixRealKCM_Freq500_uid89_T1_Freq500_uid95
-- VHDL generated for DummyFPGA @ 500MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 2
-- Target frequency (MHz): 500
-- Input signals: X
-- Output signals: Y
--  approx. input signal timings: X: (c0, 0.000000ns)
--  approx. output signal timings: Y: (c0, 0.550000ns)

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity FixRealKCM_Freq500_uid89_T1_Freq500_uid95 is
    port (X : in  std_logic_vector(2 downto 0);
          Y : out  std_logic_vector(12 downto 0)   );
end entity;

architecture arch of FixRealKCM_Freq500_uid89_T1_Freq500_uid95 is
signal Y0 :  std_logic_vector(12 downto 0);
   -- timing of Y0: (c0, 0.550000ns)
signal Y1 :  std_logic_vector(12 downto 0);
   -- timing of Y1: (c0, 0.550000ns)
begin
   with X  select  Y0 <= 
      "0000000000000" when "000",
      "0001011000110" when "001",
      "0010110001100" when "010",
      "0100001010001" when "011",
      "0101100010111" when "100",
      "0110111011101" when "101",
      "1000010100011" when "110",
      "1001101101000" when "111",
      "-------------" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                     FixFunctionByTable_Freq500_uid104
-- Evaluator for exp(x*1b-1) on [-1,1) for lsbIn=-9 (wIn=10), msbout=0, lsbOut=-12 (wOut=13). Out interval: [0.606531; 1.64711]. Output is unsigned

-- VHDL generated for DummyFPGA @ 500MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin (2010-2018)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 2
-- Target frequency (MHz): 500
-- Input signals: X
-- Output signals: Y
--  approx. input signal timings: X: (c0, 0.000000ns)
--  approx. output signal timings: Y: (c0, 0.550000ns)

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity FixFunctionByTable_Freq500_uid104 is
    port (X : in  std_logic_vector(9 downto 0);
          Y : out  std_logic_vector(12 downto 0)   );
end entity;

architecture arch of FixFunctionByTable_Freq500_uid104 is
signal Y0 :  std_logic_vector(12 downto 0);
   -- timing of Y0: (c0, 0.550000ns)
signal Y1 :  std_logic_vector(12 downto 0);
   -- timing of Y1: (c0, 0.550000ns)
begin
   with X  select  Y0 <= 
      "1000000000000" when "0000000000",
      "1000000000100" when "0000000001",
      "1000000001000" when "0000000010",
      "1000000001100" when "0000000011",
      "1000000010000" when "0000000100",
      "1000000010100" when "0000000101",
      "1000000011000" when "0000000110",
      "1000000011100" when "0000000111",
      "1000000100000" when "0000001000",
      "1000000100100" when "0000001001",
      "1000000101000" when "0000001010",
      "1000000101100" when "0000001011",
      "1000000110000" when "0000001100",
      "1000000110100" when "0000001101",
      "1000000111000" when "0000001110",
      "1000000111100" when "0000001111",
      "1000001000001" when "0000010000",
      "1000001000101" when "0000010001",
      "1000001001001" when "0000010010",
      "1000001001101" when "0000010011",
      "1000001010001" when "0000010100",
      "1000001010101" when "0000010101",
      "1000001011001" when "0000010110",
      "1000001011101" when "0000010111",
      "1000001100001" when "0000011000",
      "1000001100101" when "0000011001",
      "1000001101001" when "0000011010",
      "1000001101101" when "0000011011",
      "1000001110010" when "0000011100",
      "1000001110110" when "0000011101",
      "1000001111010" when "0000011110",
      "1000001111110" when "0000011111",
      "1000010000010" when "0000100000",
      "1000010000110" when "0000100001",
      "1000010001010" when "0000100010",
      "1000010001110" when "0000100011",
      "1000010010011" when "0000100100",
      "1000010010111" when "0000100101",
      "1000010011011" when "0000100110",
      "1000010011111" when "0000100111",
      "1000010100011" when "0000101000",
      "1000010100111" when "0000101001",
      "1000010101011" when "0000101010",
      "1000010110000" when "0000101011",
      "1000010110100" when "0000101100",
      "1000010111000" when "0000101101",
      "1000010111100" when "0000101110",
      "1000011000000" when "0000101111",
      "1000011000101" when "0000110000",
      "1000011001001" when "0000110001",
      "1000011001101" when "0000110010",
      "1000011010001" when "0000110011",
      "1000011010101" when "0000110100",
      "1000011011010" when "0000110101",
      "1000011011110" when "0000110110",
      "1000011100010" when "0000110111",
      "1000011100110" when "0000111000",
      "1000011101010" when "0000111001",
      "1000011101111" when "0000111010",
      "1000011110011" when "0000111011",
      "1000011110111" when "0000111100",
      "1000011111011" when "0000111101",
      "1000100000000" when "0000111110",
      "1000100000100" when "0000111111",
      "1000100001000" when "0001000000",
      "1000100001100" when "0001000001",
      "1000100010001" when "0001000010",
      "1000100010101" when "0001000011",
      "1000100011001" when "0001000100",
      "1000100011110" when "0001000101",
      "1000100100010" when "0001000110",
      "1000100100110" when "0001000111",
      "1000100101010" when "0001001000",
      "1000100101111" when "0001001001",
      "1000100110011" when "0001001010",
      "1000100110111" when "0001001011",
      "1000100111100" when "0001001100",
      "1000101000000" when "0001001101",
      "1000101000100" when "0001001110",
      "1000101001001" when "0001001111",
      "1000101001101" when "0001010000",
      "1000101010001" when "0001010001",
      "1000101010101" when "0001010010",
      "1000101011010" when "0001010011",
      "1000101011110" when "0001010100",
      "1000101100011" when "0001010101",
      "1000101100111" when "0001010110",
      "1000101101011" when "0001010111",
      "1000101110000" when "0001011000",
      "1000101110100" when "0001011001",
      "1000101111000" when "0001011010",
      "1000101111101" when "0001011011",
      "1000110000001" when "0001011100",
      "1000110000101" when "0001011101",
      "1000110001010" when "0001011110",
      "1000110001110" when "0001011111",
      "1000110010011" when "0001100000",
      "1000110010111" when "0001100001",
      "1000110011011" when "0001100010",
      "1000110100000" when "0001100011",
      "1000110100100" when "0001100100",
      "1000110101001" when "0001100101",
      "1000110101101" when "0001100110",
      "1000110110001" when "0001100111",
      "1000110110110" when "0001101000",
      "1000110111010" when "0001101001",
      "1000110111111" when "0001101010",
      "1000111000011" when "0001101011",
      "1000111001000" when "0001101100",
      "1000111001100" when "0001101101",
      "1000111010001" when "0001101110",
      "1000111010101" when "0001101111",
      "1000111011001" when "0001110000",
      "1000111011110" when "0001110001",
      "1000111100010" when "0001110010",
      "1000111100111" when "0001110011",
      "1000111101011" when "0001110100",
      "1000111110000" when "0001110101",
      "1000111110100" when "0001110110",
      "1000111111001" when "0001110111",
      "1000111111101" when "0001111000",
      "1001000000010" when "0001111001",
      "1001000000110" when "0001111010",
      "1001000001011" when "0001111011",
      "1001000001111" when "0001111100",
      "1001000010100" when "0001111101",
      "1001000011000" when "0001111110",
      "1001000011101" when "0001111111",
      "1001000100001" when "0010000000",
      "1001000100110" when "0010000001",
      "1001000101010" when "0010000010",
      "1001000101111" when "0010000011",
      "1001000110100" when "0010000100",
      "1001000111000" when "0010000101",
      "1001000111101" when "0010000110",
      "1001001000001" when "0010000111",
      "1001001000110" when "0010001000",
      "1001001001010" when "0010001001",
      "1001001001111" when "0010001010",
      "1001001010100" when "0010001011",
      "1001001011000" when "0010001100",
      "1001001011101" when "0010001101",
      "1001001100001" when "0010001110",
      "1001001100110" when "0010001111",
      "1001001101010" when "0010010000",
      "1001001101111" when "0010010001",
      "1001001110100" when "0010010010",
      "1001001111000" when "0010010011",
      "1001001111101" when "0010010100",
      "1001010000010" when "0010010101",
      "1001010000110" when "0010010110",
      "1001010001011" when "0010010111",
      "1001010001111" when "0010011000",
      "1001010010100" when "0010011001",
      "1001010011001" when "0010011010",
      "1001010011101" when "0010011011",
      "1001010100010" when "0010011100",
      "1001010100111" when "0010011101",
      "1001010101011" when "0010011110",
      "1001010110000" when "0010011111",
      "1001010110101" when "0010100000",
      "1001010111001" when "0010100001",
      "1001010111110" when "0010100010",
      "1001011000011" when "0010100011",
      "1001011000111" when "0010100100",
      "1001011001100" when "0010100101",
      "1001011010001" when "0010100110",
      "1001011010110" when "0010100111",
      "1001011011010" when "0010101000",
      "1001011011111" when "0010101001",
      "1001011100100" when "0010101010",
      "1001011101000" when "0010101011",
      "1001011101101" when "0010101100",
      "1001011110010" when "0010101101",
      "1001011110111" when "0010101110",
      "1001011111011" when "0010101111",
      "1001100000000" when "0010110000",
      "1001100000101" when "0010110001",
      "1001100001010" when "0010110010",
      "1001100001110" when "0010110011",
      "1001100010011" when "0010110100",
      "1001100011000" when "0010110101",
      "1001100011101" when "0010110110",
      "1001100100001" when "0010110111",
      "1001100100110" when "0010111000",
      "1001100101011" when "0010111001",
      "1001100110000" when "0010111010",
      "1001100110101" when "0010111011",
      "1001100111001" when "0010111100",
      "1001100111110" when "0010111101",
      "1001101000011" when "0010111110",
      "1001101001000" when "0010111111",
      "1001101001101" when "0011000000",
      "1001101010010" when "0011000001",
      "1001101010110" when "0011000010",
      "1001101011011" when "0011000011",
      "1001101100000" when "0011000100",
      "1001101100101" when "0011000101",
      "1001101101010" when "0011000110",
      "1001101101111" when "0011000111",
      "1001101110011" when "0011001000",
      "1001101111000" when "0011001001",
      "1001101111101" when "0011001010",
      "1001110000010" when "0011001011",
      "1001110000111" when "0011001100",
      "1001110001100" when "0011001101",
      "1001110010001" when "0011001110",
      "1001110010110" when "0011001111",
      "1001110011011" when "0011010000",
      "1001110011111" when "0011010001",
      "1001110100100" when "0011010010",
      "1001110101001" when "0011010011",
      "1001110101110" when "0011010100",
      "1001110110011" when "0011010101",
      "1001110111000" when "0011010110",
      "1001110111101" when "0011010111",
      "1001111000010" when "0011011000",
      "1001111000111" when "0011011001",
      "1001111001100" when "0011011010",
      "1001111010001" when "0011011011",
      "1001111010110" when "0011011100",
      "1001111011011" when "0011011101",
      "1001111100000" when "0011011110",
      "1001111100101" when "0011011111",
      "1001111101010" when "0011100000",
      "1001111101111" when "0011100001",
      "1001111110100" when "0011100010",
      "1001111111001" when "0011100011",
      "1001111111110" when "0011100100",
      "1010000000011" when "0011100101",
      "1010000001000" when "0011100110",
      "1010000001101" when "0011100111",
      "1010000010010" when "0011101000",
      "1010000010111" when "0011101001",
      "1010000011100" when "0011101010",
      "1010000100001" when "0011101011",
      "1010000100110" when "0011101100",
      "1010000101011" when "0011101101",
      "1010000110000" when "0011101110",
      "1010000110101" when "0011101111",
      "1010000111010" when "0011110000",
      "1010000111111" when "0011110001",
      "1010001000100" when "0011110010",
      "1010001001001" when "0011110011",
      "1010001001110" when "0011110100",
      "1010001010011" when "0011110101",
      "1010001011000" when "0011110110",
      "1010001011101" when "0011110111",
      "1010001100010" when "0011111000",
      "1010001101000" when "0011111001",
      "1010001101101" when "0011111010",
      "1010001110010" when "0011111011",
      "1010001110111" when "0011111100",
      "1010001111100" when "0011111101",
      "1010010000001" when "0011111110",
      "1010010000110" when "0011111111",
      "1010010001011" when "0100000000",
      "1010010010001" when "0100000001",
      "1010010010110" when "0100000010",
      "1010010011011" when "0100000011",
      "1010010100000" when "0100000100",
      "1010010100101" when "0100000101",
      "1010010101010" when "0100000110",
      "1010010101111" when "0100000111",
      "1010010110101" when "0100001000",
      "1010010111010" when "0100001001",
      "1010010111111" when "0100001010",
      "1010011000100" when "0100001011",
      "1010011001001" when "0100001100",
      "1010011001111" when "0100001101",
      "1010011010100" when "0100001110",
      "1010011011001" when "0100001111",
      "1010011011110" when "0100010000",
      "1010011100011" when "0100010001",
      "1010011101001" when "0100010010",
      "1010011101110" when "0100010011",
      "1010011110011" when "0100010100",
      "1010011111000" when "0100010101",
      "1010011111110" when "0100010110",
      "1010100000011" when "0100010111",
      "1010100001000" when "0100011000",
      "1010100001101" when "0100011001",
      "1010100010011" when "0100011010",
      "1010100011000" when "0100011011",
      "1010100011101" when "0100011100",
      "1010100100010" when "0100011101",
      "1010100101000" when "0100011110",
      "1010100101101" when "0100011111",
      "1010100110010" when "0100100000",
      "1010100111000" when "0100100001",
      "1010100111101" when "0100100010",
      "1010101000010" when "0100100011",
      "1010101001000" when "0100100100",
      "1010101001101" when "0100100101",
      "1010101010010" when "0100100110",
      "1010101011000" when "0100100111",
      "1010101011101" when "0100101000",
      "1010101100010" when "0100101001",
      "1010101101000" when "0100101010",
      "1010101101101" when "0100101011",
      "1010101110010" when "0100101100",
      "1010101111000" when "0100101101",
      "1010101111101" when "0100101110",
      "1010110000010" when "0100101111",
      "1010110001000" when "0100110000",
      "1010110001101" when "0100110001",
      "1010110010011" when "0100110010",
      "1010110011000" when "0100110011",
      "1010110011101" when "0100110100",
      "1010110100011" when "0100110101",
      "1010110101000" when "0100110110",
      "1010110101110" when "0100110111",
      "1010110110011" when "0100111000",
      "1010110111000" when "0100111001",
      "1010110111110" when "0100111010",
      "1010111000011" when "0100111011",
      "1010111001001" when "0100111100",
      "1010111001110" when "0100111101",
      "1010111010100" when "0100111110",
      "1010111011001" when "0100111111",
      "1010111011111" when "0101000000",
      "1010111100100" when "0101000001",
      "1010111101010" when "0101000010",
      "1010111101111" when "0101000011",
      "1010111110100" when "0101000100",
      "1010111111010" when "0101000101",
      "1010111111111" when "0101000110",
      "1011000000101" when "0101000111",
      "1011000001010" when "0101001000",
      "1011000010000" when "0101001001",
      "1011000010110" when "0101001010",
      "1011000011011" when "0101001011",
      "1011000100001" when "0101001100",
      "1011000100110" when "0101001101",
      "1011000101100" when "0101001110",
      "1011000110001" when "0101001111",
      "1011000110111" when "0101010000",
      "1011000111100" when "0101010001",
      "1011001000010" when "0101010010",
      "1011001000111" when "0101010011",
      "1011001001101" when "0101010100",
      "1011001010011" when "0101010101",
      "1011001011000" when "0101010110",
      "1011001011110" when "0101010111",
      "1011001100011" when "0101011000",
      "1011001101001" when "0101011001",
      "1011001101111" when "0101011010",
      "1011001110100" when "0101011011",
      "1011001111010" when "0101011100",
      "1011001111111" when "0101011101",
      "1011010000101" when "0101011110",
      "1011010001011" when "0101011111",
      "1011010010000" when "0101100000",
      "1011010010110" when "0101100001",
      "1011010011100" when "0101100010",
      "1011010100001" when "0101100011",
      "1011010100111" when "0101100100",
      "1011010101101" when "0101100101",
      "1011010110010" when "0101100110",
      "1011010111000" when "0101100111",
      "1011010111110" when "0101101000",
      "1011011000011" when "0101101001",
      "1011011001001" when "0101101010",
      "1011011001111" when "0101101011",
      "1011011010100" when "0101101100",
      "1011011011010" when "0101101101",
      "1011011100000" when "0101101110",
      "1011011100110" when "0101101111",
      "1011011101011" when "0101110000",
      "1011011110001" when "0101110001",
      "1011011110111" when "0101110010",
      "1011011111100" when "0101110011",
      "1011100000010" when "0101110100",
      "1011100001000" when "0101110101",
      "1011100001110" when "0101110110",
      "1011100010011" when "0101110111",
      "1011100011001" when "0101111000",
      "1011100011111" when "0101111001",
      "1011100100101" when "0101111010",
      "1011100101011" when "0101111011",
      "1011100110000" when "0101111100",
      "1011100110110" when "0101111101",
      "1011100111100" when "0101111110",
      "1011101000010" when "0101111111",
      "1011101001000" when "0110000000",
      "1011101001101" when "0110000001",
      "1011101010011" when "0110000010",
      "1011101011001" when "0110000011",
      "1011101011111" when "0110000100",
      "1011101100101" when "0110000101",
      "1011101101011" when "0110000110",
      "1011101110001" when "0110000111",
      "1011101110110" when "0110001000",
      "1011101111100" when "0110001001",
      "1011110000010" when "0110001010",
      "1011110001000" when "0110001011",
      "1011110001110" when "0110001100",
      "1011110010100" when "0110001101",
      "1011110011010" when "0110001110",
      "1011110100000" when "0110001111",
      "1011110100101" when "0110010000",
      "1011110101011" when "0110010001",
      "1011110110001" when "0110010010",
      "1011110110111" when "0110010011",
      "1011110111101" when "0110010100",
      "1011111000011" when "0110010101",
      "1011111001001" when "0110010110",
      "1011111001111" when "0110010111",
      "1011111010101" when "0110011000",
      "1011111011011" when "0110011001",
      "1011111100001" when "0110011010",
      "1011111100111" when "0110011011",
      "1011111101101" when "0110011100",
      "1011111110011" when "0110011101",
      "1011111111001" when "0110011110",
      "1011111111111" when "0110011111",
      "1100000000101" when "0110100000",
      "1100000001011" when "0110100001",
      "1100000010001" when "0110100010",
      "1100000010111" when "0110100011",
      "1100000011101" when "0110100100",
      "1100000100011" when "0110100101",
      "1100000101001" when "0110100110",
      "1100000101111" when "0110100111",
      "1100000110101" when "0110101000",
      "1100000111011" when "0110101001",
      "1100001000001" when "0110101010",
      "1100001000111" when "0110101011",
      "1100001001101" when "0110101100",
      "1100001010011" when "0110101101",
      "1100001011001" when "0110101110",
      "1100001100000" when "0110101111",
      "1100001100110" when "0110110000",
      "1100001101100" when "0110110001",
      "1100001110010" when "0110110010",
      "1100001111000" when "0110110011",
      "1100001111110" when "0110110100",
      "1100010000100" when "0110110101",
      "1100010001010" when "0110110110",
      "1100010010000" when "0110110111",
      "1100010010111" when "0110111000",
      "1100010011101" when "0110111001",
      "1100010100011" when "0110111010",
      "1100010101001" when "0110111011",
      "1100010101111" when "0110111100",
      "1100010110101" when "0110111101",
      "1100010111100" when "0110111110",
      "1100011000010" when "0110111111",
      "1100011001000" when "0111000000",
      "1100011001110" when "0111000001",
      "1100011010100" when "0111000010",
      "1100011011011" when "0111000011",
      "1100011100001" when "0111000100",
      "1100011100111" when "0111000101",
      "1100011101101" when "0111000110",
      "1100011110100" when "0111000111",
      "1100011111010" when "0111001000",
      "1100100000000" when "0111001001",
      "1100100000110" when "0111001010",
      "1100100001101" when "0111001011",
      "1100100010011" when "0111001100",
      "1100100011001" when "0111001101",
      "1100100011111" when "0111001110",
      "1100100100110" when "0111001111",
      "1100100101100" when "0111010000",
      "1100100110010" when "0111010001",
      "1100100111001" when "0111010010",
      "1100100111111" when "0111010011",
      "1100101000101" when "0111010100",
      "1100101001011" when "0111010101",
      "1100101010010" when "0111010110",
      "1100101011000" when "0111010111",
      "1100101011110" when "0111011000",
      "1100101100101" when "0111011001",
      "1100101101011" when "0111011010",
      "1100101110010" when "0111011011",
      "1100101111000" when "0111011100",
      "1100101111110" when "0111011101",
      "1100110000101" when "0111011110",
      "1100110001011" when "0111011111",
      "1100110010001" when "0111100000",
      "1100110011000" when "0111100001",
      "1100110011110" when "0111100010",
      "1100110100101" when "0111100011",
      "1100110101011" when "0111100100",
      "1100110110001" when "0111100101",
      "1100110111000" when "0111100110",
      "1100110111110" when "0111100111",
      "1100111000101" when "0111101000",
      "1100111001011" when "0111101001",
      "1100111010010" when "0111101010",
      "1100111011000" when "0111101011",
      "1100111011111" when "0111101100",
      "1100111100101" when "0111101101",
      "1100111101011" when "0111101110",
      "1100111110010" when "0111101111",
      "1100111111000" when "0111110000",
      "1100111111111" when "0111110001",
      "1101000000101" when "0111110010",
      "1101000001100" when "0111110011",
      "1101000010010" when "0111110100",
      "1101000011001" when "0111110101",
      "1101000100000" when "0111110110",
      "1101000100110" when "0111110111",
      "1101000101101" when "0111111000",
      "1101000110011" when "0111111001",
      "1101000111010" when "0111111010",
      "1101001000000" when "0111111011",
      "1101001000111" when "0111111100",
      "1101001001101" when "0111111101",
      "1101001010100" when "0111111110",
      "1101001011011" when "0111111111",
      "0100110110100" when "1000000000",
      "0100110110111" when "1000000001",
      "0100110111001" when "1000000010",
      "0100110111100" when "1000000011",
      "0100110111110" when "1000000100",
      "0100111000001" when "1000000101",
      "0100111000011" when "1000000110",
      "0100111000101" when "1000000111",
      "0100111001000" when "1000001000",
      "0100111001010" when "1000001001",
      "0100111001101" when "1000001010",
      "0100111001111" when "1000001011",
      "0100111010010" when "1000001100",
      "0100111010100" when "1000001101",
      "0100111010111" when "1000001110",
      "0100111011001" when "1000001111",
      "0100111011011" when "1000010000",
      "0100111011110" when "1000010001",
      "0100111100000" when "1000010010",
      "0100111100011" when "1000010011",
      "0100111100101" when "1000010100",
      "0100111101000" when "1000010101",
      "0100111101010" when "1000010110",
      "0100111101101" when "1000010111",
      "0100111101111" when "1000011000",
      "0100111110010" when "1000011001",
      "0100111110100" when "1000011010",
      "0100111110111" when "1000011011",
      "0100111111001" when "1000011100",
      "0100111111100" when "1000011101",
      "0100111111110" when "1000011110",
      "0101000000001" when "1000011111",
      "0101000000011" when "1000100000",
      "0101000000110" when "1000100001",
      "0101000001000" when "1000100010",
      "0101000001011" when "1000100011",
      "0101000001101" when "1000100100",
      "0101000010000" when "1000100101",
      "0101000010010" when "1000100110",
      "0101000010101" when "1000100111",
      "0101000010111" when "1000101000",
      "0101000011010" when "1000101001",
      "0101000011100" when "1000101010",
      "0101000011111" when "1000101011",
      "0101000100001" when "1000101100",
      "0101000100100" when "1000101101",
      "0101000100110" when "1000101110",
      "0101000101001" when "1000101111",
      "0101000101100" when "1000110000",
      "0101000101110" when "1000110001",
      "0101000110001" when "1000110010",
      "0101000110011" when "1000110011",
      "0101000110110" when "1000110100",
      "0101000111000" when "1000110101",
      "0101000111011" when "1000110110",
      "0101000111101" when "1000110111",
      "0101001000000" when "1000111000",
      "0101001000011" when "1000111001",
      "0101001000101" when "1000111010",
      "0101001001000" when "1000111011",
      "0101001001010" when "1000111100",
      "0101001001101" when "1000111101",
      "0101001001111" when "1000111110",
      "0101001010010" when "1000111111",
      "0101001010101" when "1001000000",
      "0101001010111" when "1001000001",
      "0101001011010" when "1001000010",
      "0101001011100" when "1001000011",
      "0101001011111" when "1001000100",
      "0101001100010" when "1001000101",
      "0101001100100" when "1001000110",
      "0101001100111" when "1001000111",
      "0101001101001" when "1001001000",
      "0101001101100" when "1001001001",
      "0101001101111" when "1001001010",
      "0101001110001" when "1001001011",
      "0101001110100" when "1001001100",
      "0101001110110" when "1001001101",
      "0101001111001" when "1001001110",
      "0101001111100" when "1001001111",
      "0101001111110" when "1001010000",
      "0101010000001" when "1001010001",
      "0101010000011" when "1001010010",
      "0101010000110" when "1001010011",
      "0101010001001" when "1001010100",
      "0101010001011" when "1001010101",
      "0101010001110" when "1001010110",
      "0101010010001" when "1001010111",
      "0101010010011" when "1001011000",
      "0101010010110" when "1001011001",
      "0101010011001" when "1001011010",
      "0101010011011" when "1001011011",
      "0101010011110" when "1001011100",
      "0101010100001" when "1001011101",
      "0101010100011" when "1001011110",
      "0101010100110" when "1001011111",
      "0101010101001" when "1001100000",
      "0101010101011" when "1001100001",
      "0101010101110" when "1001100010",
      "0101010110001" when "1001100011",
      "0101010110011" when "1001100100",
      "0101010110110" when "1001100101",
      "0101010111001" when "1001100110",
      "0101010111011" when "1001100111",
      "0101010111110" when "1001101000",
      "0101011000001" when "1001101001",
      "0101011000011" when "1001101010",
      "0101011000110" when "1001101011",
      "0101011001001" when "1001101100",
      "0101011001011" when "1001101101",
      "0101011001110" when "1001101110",
      "0101011010001" when "1001101111",
      "0101011010011" when "1001110000",
      "0101011010110" when "1001110001",
      "0101011011001" when "1001110010",
      "0101011011100" when "1001110011",
      "0101011011110" when "1001110100",
      "0101011100001" when "1001110101",
      "0101011100100" when "1001110110",
      "0101011100111" when "1001110111",
      "0101011101001" when "1001111000",
      "0101011101100" when "1001111001",
      "0101011101111" when "1001111010",
      "0101011110001" when "1001111011",
      "0101011110100" when "1001111100",
      "0101011110111" when "1001111101",
      "0101011111010" when "1001111110",
      "0101011111100" when "1001111111",
      "0101011111111" when "1010000000",
      "0101100000010" when "1010000001",
      "0101100000101" when "1010000010",
      "0101100000111" when "1010000011",
      "0101100001010" when "1010000100",
      "0101100001101" when "1010000101",
      "0101100010000" when "1010000110",
      "0101100010010" when "1010000111",
      "0101100010101" when "1010001000",
      "0101100011000" when "1010001001",
      "0101100011011" when "1010001010",
      "0101100011110" when "1010001011",
      "0101100100000" when "1010001100",
      "0101100100011" when "1010001101",
      "0101100100110" when "1010001110",
      "0101100101001" when "1010001111",
      "0101100101011" when "1010010000",
      "0101100101110" when "1010010001",
      "0101100110001" when "1010010010",
      "0101100110100" when "1010010011",
      "0101100110111" when "1010010100",
      "0101100111001" when "1010010101",
      "0101100111100" when "1010010110",
      "0101100111111" when "1010010111",
      "0101101000010" when "1010011000",
      "0101101000101" when "1010011001",
      "0101101001000" when "1010011010",
      "0101101001010" when "1010011011",
      "0101101001101" when "1010011100",
      "0101101010000" when "1010011101",
      "0101101010011" when "1010011110",
      "0101101010110" when "1010011111",
      "0101101011000" when "1010100000",
      "0101101011011" when "1010100001",
      "0101101011110" when "1010100010",
      "0101101100001" when "1010100011",
      "0101101100100" when "1010100100",
      "0101101100111" when "1010100101",
      "0101101101010" when "1010100110",
      "0101101101100" when "1010100111",
      "0101101101111" when "1010101000",
      "0101101110010" when "1010101001",
      "0101101110101" when "1010101010",
      "0101101111000" when "1010101011",
      "0101101111011" when "1010101100",
      "0101101111110" when "1010101101",
      "0101110000000" when "1010101110",
      "0101110000011" when "1010101111",
      "0101110000110" when "1010110000",
      "0101110001001" when "1010110001",
      "0101110001100" when "1010110010",
      "0101110001111" when "1010110011",
      "0101110010010" when "1010110100",
      "0101110010101" when "1010110101",
      "0101110011000" when "1010110110",
      "0101110011010" when "1010110111",
      "0101110011101" when "1010111000",
      "0101110100000" when "1010111001",
      "0101110100011" when "1010111010",
      "0101110100110" when "1010111011",
      "0101110101001" when "1010111100",
      "0101110101100" when "1010111101",
      "0101110101111" when "1010111110",
      "0101110110010" when "1010111111",
      "0101110110101" when "1011000000",
      "0101110111000" when "1011000001",
      "0101110111011" when "1011000010",
      "0101110111101" when "1011000011",
      "0101111000000" when "1011000100",
      "0101111000011" when "1011000101",
      "0101111000110" when "1011000110",
      "0101111001001" when "1011000111",
      "0101111001100" when "1011001000",
      "0101111001111" when "1011001001",
      "0101111010010" when "1011001010",
      "0101111010101" when "1011001011",
      "0101111011000" when "1011001100",
      "0101111011011" when "1011001101",
      "0101111011110" when "1011001110",
      "0101111100001" when "1011001111",
      "0101111100100" when "1011010000",
      "0101111100111" when "1011010001",
      "0101111101010" when "1011010010",
      "0101111101101" when "1011010011",
      "0101111110000" when "1011010100",
      "0101111110011" when "1011010101",
      "0101111110110" when "1011010110",
      "0101111111001" when "1011010111",
      "0101111111100" when "1011011000",
      "0101111111111" when "1011011001",
      "0110000000010" when "1011011010",
      "0110000000101" when "1011011011",
      "0110000001000" when "1011011100",
      "0110000001011" when "1011011101",
      "0110000001110" when "1011011110",
      "0110000010001" when "1011011111",
      "0110000010100" when "1011100000",
      "0110000010111" when "1011100001",
      "0110000011010" when "1011100010",
      "0110000011101" when "1011100011",
      "0110000100000" when "1011100100",
      "0110000100011" when "1011100101",
      "0110000100110" when "1011100110",
      "0110000101001" when "1011100111",
      "0110000101100" when "1011101000",
      "0110000101111" when "1011101001",
      "0110000110010" when "1011101010",
      "0110000110101" when "1011101011",
      "0110000111000" when "1011101100",
      "0110000111011" when "1011101101",
      "0110000111110" when "1011101110",
      "0110001000001" when "1011101111",
      "0110001000101" when "1011110000",
      "0110001001000" when "1011110001",
      "0110001001011" when "1011110010",
      "0110001001110" when "1011110011",
      "0110001010001" when "1011110100",
      "0110001010100" when "1011110101",
      "0110001010111" when "1011110110",
      "0110001011010" when "1011110111",
      "0110001011101" when "1011111000",
      "0110001100000" when "1011111001",
      "0110001100011" when "1011111010",
      "0110001100110" when "1011111011",
      "0110001101010" when "1011111100",
      "0110001101101" when "1011111101",
      "0110001110000" when "1011111110",
      "0110001110011" when "1011111111",
      "0110001110110" when "1100000000",
      "0110001111001" when "1100000001",
      "0110001111100" when "1100000010",
      "0110001111111" when "1100000011",
      "0110010000010" when "1100000100",
      "0110010000110" when "1100000101",
      "0110010001001" when "1100000110",
      "0110010001100" when "1100000111",
      "0110010001111" when "1100001000",
      "0110010010010" when "1100001001",
      "0110010010101" when "1100001010",
      "0110010011000" when "1100001011",
      "0110010011100" when "1100001100",
      "0110010011111" when "1100001101",
      "0110010100010" when "1100001110",
      "0110010100101" when "1100001111",
      "0110010101000" when "1100010000",
      "0110010101011" when "1100010001",
      "0110010101111" when "1100010010",
      "0110010110010" when "1100010011",
      "0110010110101" when "1100010100",
      "0110010111000" when "1100010101",
      "0110010111011" when "1100010110",
      "0110010111110" when "1100010111",
      "0110011000010" when "1100011000",
      "0110011000101" when "1100011001",
      "0110011001000" when "1100011010",
      "0110011001011" when "1100011011",
      "0110011001110" when "1100011100",
      "0110011010010" when "1100011101",
      "0110011010101" when "1100011110",
      "0110011011000" when "1100011111",
      "0110011011011" when "1100100000",
      "0110011011110" when "1100100001",
      "0110011100010" when "1100100010",
      "0110011100101" when "1100100011",
      "0110011101000" when "1100100100",
      "0110011101011" when "1100100101",
      "0110011101111" when "1100100110",
      "0110011110010" when "1100100111",
      "0110011110101" when "1100101000",
      "0110011111000" when "1100101001",
      "0110011111100" when "1100101010",
      "0110011111111" when "1100101011",
      "0110100000010" when "1100101100",
      "0110100000101" when "1100101101",
      "0110100001001" when "1100101110",
      "0110100001100" when "1100101111",
      "0110100001111" when "1100110000",
      "0110100010010" when "1100110001",
      "0110100010110" when "1100110010",
      "0110100011001" when "1100110011",
      "0110100011100" when "1100110100",
      "0110100011111" when "1100110101",
      "0110100100011" when "1100110110",
      "0110100100110" when "1100110111",
      "0110100101001" when "1100111000",
      "0110100101101" when "1100111001",
      "0110100110000" when "1100111010",
      "0110100110011" when "1100111011",
      "0110100110110" when "1100111100",
      "0110100111010" when "1100111101",
      "0110100111101" when "1100111110",
      "0110101000000" when "1100111111",
      "0110101000100" when "1101000000",
      "0110101000111" when "1101000001",
      "0110101001010" when "1101000010",
      "0110101001110" when "1101000011",
      "0110101010001" when "1101000100",
      "0110101010100" when "1101000101",
      "0110101011000" when "1101000110",
      "0110101011011" when "1101000111",
      "0110101011110" when "1101001000",
      "0110101100010" when "1101001001",
      "0110101100101" when "1101001010",
      "0110101101000" when "1101001011",
      "0110101101100" when "1101001100",
      "0110101101111" when "1101001101",
      "0110101110010" when "1101001110",
      "0110101110110" when "1101001111",
      "0110101111001" when "1101010000",
      "0110101111101" when "1101010001",
      "0110110000000" when "1101010010",
      "0110110000011" when "1101010011",
      "0110110000111" when "1101010100",
      "0110110001010" when "1101010101",
      "0110110001101" when "1101010110",
      "0110110010001" when "1101010111",
      "0110110010100" when "1101011000",
      "0110110011000" when "1101011001",
      "0110110011011" when "1101011010",
      "0110110011110" when "1101011011",
      "0110110100010" when "1101011100",
      "0110110100101" when "1101011101",
      "0110110101001" when "1101011110",
      "0110110101100" when "1101011111",
      "0110110101111" when "1101100000",
      "0110110110011" when "1101100001",
      "0110110110110" when "1101100010",
      "0110110111010" when "1101100011",
      "0110110111101" when "1101100100",
      "0110111000001" when "1101100101",
      "0110111000100" when "1101100110",
      "0110111001000" when "1101100111",
      "0110111001011" when "1101101000",
      "0110111001110" when "1101101001",
      "0110111010010" when "1101101010",
      "0110111010101" when "1101101011",
      "0110111011001" when "1101101100",
      "0110111011100" when "1101101101",
      "0110111100000" when "1101101110",
      "0110111100011" when "1101101111",
      "0110111100111" when "1101110000",
      "0110111101010" when "1101110001",
      "0110111101110" when "1101110010",
      "0110111110001" when "1101110011",
      "0110111110101" when "1101110100",
      "0110111111000" when "1101110101",
      "0110111111100" when "1101110110",
      "0110111111111" when "1101110111",
      "0111000000011" when "1101111000",
      "0111000000110" when "1101111001",
      "0111000001010" when "1101111010",
      "0111000001101" when "1101111011",
      "0111000010001" when "1101111100",
      "0111000010100" when "1101111101",
      "0111000011000" when "1101111110",
      "0111000011011" when "1101111111",
      "0111000011111" when "1110000000",
      "0111000100010" when "1110000001",
      "0111000100110" when "1110000010",
      "0111000101001" when "1110000011",
      "0111000101101" when "1110000100",
      "0111000110000" when "1110000101",
      "0111000110100" when "1110000110",
      "0111000111000" when "1110000111",
      "0111000111011" when "1110001000",
      "0111000111111" when "1110001001",
      "0111001000010" when "1110001010",
      "0111001000110" when "1110001011",
      "0111001001001" when "1110001100",
      "0111001001101" when "1110001101",
      "0111001010000" when "1110001110",
      "0111001010100" when "1110001111",
      "0111001011000" when "1110010000",
      "0111001011011" when "1110010001",
      "0111001011111" when "1110010010",
      "0111001100010" when "1110010011",
      "0111001100110" when "1110010100",
      "0111001101010" when "1110010101",
      "0111001101101" when "1110010110",
      "0111001110001" when "1110010111",
      "0111001110100" when "1110011000",
      "0111001111000" when "1110011001",
      "0111001111100" when "1110011010",
      "0111001111111" when "1110011011",
      "0111010000011" when "1110011100",
      "0111010000111" when "1110011101",
      "0111010001010" when "1110011110",
      "0111010001110" when "1110011111",
      "0111010010001" when "1110100000",
      "0111010010101" when "1110100001",
      "0111010011001" when "1110100010",
      "0111010011100" when "1110100011",
      "0111010100000" when "1110100100",
      "0111010100100" when "1110100101",
      "0111010100111" when "1110100110",
      "0111010101011" when "1110100111",
      "0111010101111" when "1110101000",
      "0111010110010" when "1110101001",
      "0111010110110" when "1110101010",
      "0111010111010" when "1110101011",
      "0111010111101" when "1110101100",
      "0111011000001" when "1110101101",
      "0111011000101" when "1110101110",
      "0111011001000" when "1110101111",
      "0111011001100" when "1110110000",
      "0111011010000" when "1110110001",
      "0111011010100" when "1110110010",
      "0111011010111" when "1110110011",
      "0111011011011" when "1110110100",
      "0111011011111" when "1110110101",
      "0111011100010" when "1110110110",
      "0111011100110" when "1110110111",
      "0111011101010" when "1110111000",
      "0111011101110" when "1110111001",
      "0111011110001" when "1110111010",
      "0111011110101" when "1110111011",
      "0111011111001" when "1110111100",
      "0111011111101" when "1110111101",
      "0111100000000" when "1110111110",
      "0111100000100" when "1110111111",
      "0111100001000" when "1111000000",
      "0111100001100" when "1111000001",
      "0111100001111" when "1111000010",
      "0111100010011" when "1111000011",
      "0111100010111" when "1111000100",
      "0111100011011" when "1111000101",
      "0111100011110" when "1111000110",
      "0111100100010" when "1111000111",
      "0111100100110" when "1111001000",
      "0111100101010" when "1111001001",
      "0111100101110" when "1111001010",
      "0111100110001" when "1111001011",
      "0111100110101" when "1111001100",
      "0111100111001" when "1111001101",
      "0111100111101" when "1111001110",
      "0111101000001" when "1111001111",
      "0111101000100" when "1111010000",
      "0111101001000" when "1111010001",
      "0111101001100" when "1111010010",
      "0111101010000" when "1111010011",
      "0111101010100" when "1111010100",
      "0111101011000" when "1111010101",
      "0111101011011" when "1111010110",
      "0111101011111" when "1111010111",
      "0111101100011" when "1111011000",
      "0111101100111" when "1111011001",
      "0111101101011" when "1111011010",
      "0111101101111" when "1111011011",
      "0111101110011" when "1111011100",
      "0111101110110" when "1111011101",
      "0111101111010" when "1111011110",
      "0111101111110" when "1111011111",
      "0111110000010" when "1111100000",
      "0111110000110" when "1111100001",
      "0111110001010" when "1111100010",
      "0111110001110" when "1111100011",
      "0111110010010" when "1111100100",
      "0111110010101" when "1111100101",
      "0111110011001" when "1111100110",
      "0111110011101" when "1111100111",
      "0111110100001" when "1111101000",
      "0111110100101" when "1111101001",
      "0111110101001" when "1111101010",
      "0111110101101" when "1111101011",
      "0111110110001" when "1111101100",
      "0111110110101" when "1111101101",
      "0111110111001" when "1111101110",
      "0111110111101" when "1111101111",
      "0111111000000" when "1111110000",
      "0111111000100" when "1111110001",
      "0111111001000" when "1111110010",
      "0111111001100" when "1111110011",
      "0111111010000" when "1111110100",
      "0111111010100" when "1111110101",
      "0111111011000" when "1111110110",
      "0111111011100" when "1111110111",
      "0111111100000" when "1111111000",
      "0111111100100" when "1111111001",
      "0111111101000" when "1111111010",
      "0111111101100" when "1111111011",
      "0111111110000" when "1111111100",
      "0111111110100" when "1111111101",
      "0111111111000" when "1111111110",
      "0111111111100" when "1111111111",
      "-------------" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          IntAdder_16_Freq500_uid5
-- VHDL generated for DummyFPGA @ 500MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin (2008-2016)
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 2
-- Target frequency (MHz): 500
-- Input signals: X Y Cin
-- Output signals: R
--  approx. input signal timings: X: (c0, 0.000000ns)Y: (c0, 0.000000ns)Cin: (c0, 0.000000ns)
--  approx. output signal timings: R: (c0, 1.150000ns)

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntAdder_16_Freq500_uid5 is
    port (clk : in std_logic;
          X : in  std_logic_vector(15 downto 0);
          Y : in  std_logic_vector(15 downto 0);
          Cin : in  std_logic;
          R : out  std_logic_vector(15 downto 0)   );
end entity;

architecture arch of IntAdder_16_Freq500_uid5 is
signal Rtmp :  std_logic_vector(15 downto 0);
   -- timing of Rtmp: (c0, 1.150000ns)
begin
   Rtmp <= X + Y + Cin;
   R <= Rtmp;
end architecture;

--------------------------------------------------------------------------------
--                             LZC_7_Freq500_uid7
-- VHDL generated for DummyFPGA @ 500MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007)
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 2
-- Target frequency (MHz): 500
-- Input signals: I
-- Output signals: O
--  approx. input signal timings: I: (c0, 0.000000ns)
--  approx. output signal timings: O: (c0, 1.660000ns)

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity LZC_7_Freq500_uid7 is
    port (clk : in std_logic;
          I : in  std_logic_vector(6 downto 0);
          O : out  std_logic_vector(2 downto 0)   );
end entity;

architecture arch of LZC_7_Freq500_uid7 is
signal level3 :  std_logic_vector(6 downto 0);
   -- timing of level3: (c0, 0.000000ns)
signal digit2 :  std_logic;
   -- timing of digit2: (c0, 0.560000ns)
signal level2 :  std_logic_vector(2 downto 0);
   -- timing of level2: (c0, 1.110000ns)
signal lowBits :  std_logic_vector(1 downto 0);
   -- timing of lowBits: (c0, 1.660000ns)
signal outHighBits :  std_logic_vector(0 downto 0);
   -- timing of outHighBits: (c0, 0.560000ns)
begin
   -- pad input to the next power of two minus 1
   level3 <= I;
   -- Main iteration for large inputs
   digit2<= '1' when level3(6 downto 3) = "0000" else '0';
   level2<= level3(2 downto 0) when digit2='1' else level3(6 downto 4);
   -- Finish counting with one LUT
   with level2  select  lowBits <= 
      "11" when "000",
      "10" when "001",
      "01" when "010",
      "01" when "011",
      "00" when others;
   outHighBits <= digit2 & "";
   O <= outHighBits & lowBits ;
end architecture;

--------------------------------------------------------------------------------
--                           LZOC_17_Freq500_uid11
-- VHDL generated for DummyFPGA @ 500MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007)
--------------------------------------------------------------------------------
-- Pipeline depth: 3 cycles
-- Clock period (ns): 2
-- Target frequency (MHz): 500
-- Input signals: I OZB
-- Output signals: O
--  approx. input signal timings: I: (c0, 0.550000ns)OZB: (c0, 0.000000ns)
--  approx. output signal timings: O: (c3, 0.410000ns)

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity LZOC_17_Freq500_uid11 is
    port (clk : in std_logic;
          I : in  std_logic_vector(16 downto 0);
          OZB : in  std_logic;
          O : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of LZOC_17_Freq500_uid11 is
signal sozb, sozb_d1, sozb_d2 :  std_logic;
   -- timing of sozb: (c0, 0.000000ns)
signal level5, level5_d1 :  std_logic_vector(30 downto 0);
   -- timing of level5: (c0, 0.550000ns)
signal digit4, digit4_d1, digit4_d2 :  std_logic;
   -- timing of digit4: (c0, 1.590000ns)
signal level4, level4_d1 :  std_logic_vector(14 downto 0);
   -- timing of level4: (c1, 0.340000ns)
signal digit3, digit3_d1 :  std_logic;
   -- timing of digit3: (c1, 1.360000ns)
signal level3 :  std_logic_vector(6 downto 0);
   -- timing of level3: (c2, 0.110000ns)
signal digit2 :  std_logic;
   -- timing of digit2: (c2, 1.110000ns)
signal level2, level2_d1 :  std_logic_vector(2 downto 0);
   -- timing of level2: (c2, 1.660000ns)
signal z :  std_logic_vector(2 downto 0);
   -- timing of z: (c3, 0.410000ns)
signal lowBits :  std_logic_vector(1 downto 0);
   -- timing of lowBits: (c3, 0.410000ns)
signal outHighBits, outHighBits_d1 :  std_logic_vector(2 downto 0);
   -- timing of outHighBits: (c2, 1.110000ns)
signal OZB_d1, OZB_d2, OZB_d3 :  std_logic;
   -- timing of OZB: (c0, 0.000000ns)
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            sozb_d1 <=  sozb;
            sozb_d2 <=  sozb_d1;
            level5_d1 <=  level5;
            digit4_d1 <=  digit4;
            digit4_d2 <=  digit4_d1;
            level4_d1 <=  level4;
            digit3_d1 <=  digit3;
            level2_d1 <=  level2;
            outHighBits_d1 <=  outHighBits;
            OZB_d1 <=  OZB;
            OZB_d2 <=  OZB_d1;
            OZB_d3 <=  OZB_d2;
         end if;
      end process;
   sozb <= OZB;
   -- pad input to the next power of two minus 1
   level5 <= I & (13 downto 0 => not sozb);
   -- Main iteration for large inputs
   digit4<= '1' when level5(30 downto 15) = (15 downto 0 => sozb) else '0';
   level4<= level5_d1(14 downto 0) when digit4_d1='1' else level5_d1(30 downto 16);
   digit3<= '1' when level4(14 downto 7) = (7 downto 0 => sozb_d1) else '0';
   level3<= level4_d1(6 downto 0) when digit3_d1='1' else level4_d1(14 downto 8);
   digit2<= '1' when level3(6 downto 3) = (3 downto 0 => sozb_d2) else '0';
   level2<= level3(2 downto 0) when digit2='1' else level3(6 downto 4);
   -- Finish counting with one LUT
   z <= level2_d1 when OZB_d3='0' else (not level2_d1);
   with z  select  lowBits <= 
      "11" when "000",
      "10" when "001",
      "01" when "010",
      "01" when "011",
      "00" when others;
   outHighBits <= digit4_d2 & digit3_d1 & digit2 & "";
   O <= outHighBits_d1 & lowBits ;
end architecture;

--------------------------------------------------------------------------------
--                   LeftShifter10_by_max_10_Freq500_uid13
-- VHDL generated for DummyFPGA @ 500MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca (2008-2011), Florent de Dinechin (2008-2019)
--------------------------------------------------------------------------------
-- Pipeline depth: 4 cycles
-- Clock period (ns): 2
-- Target frequency (MHz): 500
-- Input signals: X S
-- Output signals: R
--  approx. input signal timings: X: (c0, 1.640000ns)S: (c3, 1.460000ns)
--  approx. output signal timings: R: (c4, 1.344615ns)

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity LeftShifter10_by_max_10_Freq500_uid13 is
    port (clk : in std_logic;
          X : in  std_logic_vector(9 downto 0);
          S : in  std_logic_vector(3 downto 0);
          R : out  std_logic_vector(19 downto 0)   );
end entity;

architecture arch of LeftShifter10_by_max_10_Freq500_uid13 is
signal ps, ps_d1 :  std_logic_vector(3 downto 0);
   -- timing of ps: (c3, 1.460000ns)
signal level0, level0_d1, level0_d2, level0_d3 :  std_logic_vector(9 downto 0);
   -- timing of level0: (c0, 1.640000ns)
signal level1, level1_d1 :  std_logic_vector(10 downto 0);
   -- timing of level1: (c3, 1.460000ns)
signal level2 :  std_logic_vector(12 downto 0);
   -- timing of level2: (c4, 0.410000ns)
signal level3 :  std_logic_vector(16 downto 0);
   -- timing of level3: (c4, 0.410000ns)
signal level4 :  std_logic_vector(24 downto 0);
   -- timing of level4: (c4, 1.344615ns)
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            ps_d1 <=  ps;
            level0_d1 <=  level0;
            level0_d2 <=  level0_d1;
            level0_d3 <=  level0_d2;
            level1_d1 <=  level1;
         end if;
      end process;
   ps<= S;
   level0<= X;
   level1<= level0_d3 & (0 downto 0 => '0') when ps(0)= '1' else     (0 downto 0 => '0') & level0_d3;
   level2<= level1_d1 & (1 downto 0 => '0') when ps_d1(1)= '1' else     (1 downto 0 => '0') & level1_d1;
   level3<= level2 & (3 downto 0 => '0') when ps_d1(2)= '1' else     (3 downto 0 => '0') & level2;
   level4<= level3 & (7 downto 0 => '0') when ps_d1(3)= '1' else     (7 downto 0 => '0') & level3;
   R <= level4(19 downto 0);
end architecture;

--------------------------------------------------------------------------------
--                         IntAdder_21_Freq500_uid19
-- VHDL generated for DummyFPGA @ 500MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin (2008-2016)
--------------------------------------------------------------------------------
-- Pipeline depth: 2 cycles
-- Clock period (ns): 2
-- Target frequency (MHz): 500
-- Input signals: X Y Cin
-- Output signals: R
--  approx. input signal timings: X: (c1, 0.560000ns)Y: (c1, 1.110000ns)Cin: (c0, 0.000000ns)
--  approx. output signal timings: R: (c2, 0.520000ns)

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntAdder_21_Freq500_uid19 is
    port (clk : in std_logic;
          X : in  std_logic_vector(20 downto 0);
          Y : in  std_logic_vector(20 downto 0);
          Cin : in  std_logic;
          R : out  std_logic_vector(20 downto 0)   );
end entity;

architecture arch of IntAdder_21_Freq500_uid19 is
signal Cin_1, Cin_1_d1, Cin_1_d2 :  std_logic;
   -- timing of Cin_1: (c0, 0.000000ns)
signal X_1, X_1_d1 :  std_logic_vector(21 downto 0);
   -- timing of X_1: (c1, 0.560000ns)
signal Y_1, Y_1_d1 :  std_logic_vector(21 downto 0);
   -- timing of Y_1: (c1, 1.110000ns)
signal S_1 :  std_logic_vector(21 downto 0);
   -- timing of S_1: (c2, 0.520000ns)
signal R_1 :  std_logic_vector(20 downto 0);
   -- timing of R_1: (c2, 0.520000ns)
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            Cin_1_d1 <=  Cin_1;
            Cin_1_d2 <=  Cin_1_d1;
            X_1_d1 <=  X_1;
            Y_1_d1 <=  Y_1;
         end if;
      end process;
   Cin_1 <= Cin;
   X_1 <= '0' & X(20 downto 0);
   Y_1 <= '0' & Y(20 downto 0);
   S_1 <= X_1_d1 + Y_1_d1 + Cin_1_d2;
   R_1 <= S_1(20 downto 0);
   R <= R_1 ;
end architecture;

--------------------------------------------------------------------------------
--                         IntAdder_21_Freq500_uid22
-- VHDL generated for DummyFPGA @ 500MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin (2008-2016)
--------------------------------------------------------------------------------
-- Pipeline depth: 3 cycles
-- Clock period (ns): 2
-- Target frequency (MHz): 500
-- Input signals: X Y Cin
-- Output signals: R
--  approx. input signal timings: X: (c2, 0.520000ns)Y: (c2, 1.100000ns)Cin: (c0, 0.000000ns)
--  approx. output signal timings: R: (c3, 0.510000ns)

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntAdder_21_Freq500_uid22 is
    port (clk : in std_logic;
          X : in  std_logic_vector(20 downto 0);
          Y : in  std_logic_vector(20 downto 0);
          Cin : in  std_logic;
          R : out  std_logic_vector(20 downto 0)   );
end entity;

architecture arch of IntAdder_21_Freq500_uid22 is
signal Cin_1, Cin_1_d1, Cin_1_d2, Cin_1_d3 :  std_logic;
   -- timing of Cin_1: (c0, 0.000000ns)
signal X_1, X_1_d1 :  std_logic_vector(21 downto 0);
   -- timing of X_1: (c2, 0.520000ns)
signal Y_1, Y_1_d1 :  std_logic_vector(21 downto 0);
   -- timing of Y_1: (c2, 1.100000ns)
signal S_1 :  std_logic_vector(21 downto 0);
   -- timing of S_1: (c3, 0.510000ns)
signal R_1 :  std_logic_vector(20 downto 0);
   -- timing of R_1: (c3, 0.510000ns)
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            Cin_1_d1 <=  Cin_1;
            Cin_1_d2 <=  Cin_1_d1;
            Cin_1_d3 <=  Cin_1_d2;
            X_1_d1 <=  X_1;
            Y_1_d1 <=  Y_1;
         end if;
      end process;
   Cin_1 <= Cin;
   X_1 <= '0' & X(20 downto 0);
   Y_1 <= '0' & Y(20 downto 0);
   S_1 <= X_1_d1 + Y_1_d1 + Cin_1_d3;
   R_1 <= S_1(20 downto 0);
   R <= R_1 ;
end architecture;

--------------------------------------------------------------------------------
--                         IntAdder_21_Freq500_uid25
-- VHDL generated for DummyFPGA @ 500MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin (2008-2016)
--------------------------------------------------------------------------------
-- Pipeline depth: 6 cycles
-- Clock period (ns): 2
-- Target frequency (MHz): 500
-- Input signals: X Y Cin
-- Output signals: R
--  approx. input signal timings: X: (c3, 0.510000ns)Y: (c5, 0.644615ns)Cin: (c0, 0.000000ns)
--  approx. output signal timings: R: (c6, 0.044615ns)

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntAdder_21_Freq500_uid25 is
    port (clk : in std_logic;
          X : in  std_logic_vector(20 downto 0);
          Y : in  std_logic_vector(20 downto 0);
          Cin : in  std_logic;
          R : out  std_logic_vector(20 downto 0)   );
end entity;

architecture arch of IntAdder_21_Freq500_uid25 is
signal Rtmp :  std_logic_vector(20 downto 0);
   -- timing of Rtmp: (c6, 0.044615ns)
signal X_d1, X_d2, X_d3 :  std_logic_vector(20 downto 0);
   -- timing of X: (c3, 0.510000ns)
signal Y_d1 :  std_logic_vector(20 downto 0);
   -- timing of Y: (c5, 0.644615ns)
signal Cin_d1, Cin_d2, Cin_d3, Cin_d4, Cin_d5, Cin_d6 :  std_logic;
   -- timing of Cin: (c0, 0.000000ns)
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            X_d1 <=  X;
            X_d2 <=  X_d1;
            X_d3 <=  X_d2;
            Y_d1 <=  Y;
            Cin_d1 <=  Cin;
            Cin_d2 <=  Cin_d1;
            Cin_d3 <=  Cin_d2;
            Cin_d4 <=  Cin_d3;
            Cin_d5 <=  Cin_d4;
            Cin_d6 <=  Cin_d5;
         end if;
      end process;
   Rtmp <= X_d3 + Y_d1 + Cin_d6;
   R <= Rtmp;
end architecture;

--------------------------------------------------------------------------------
--                         IntAdder_30_Freq500_uid34
-- VHDL generated for DummyFPGA @ 500MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin (2008-2016)
--------------------------------------------------------------------------------
-- Pipeline depth: 2 cycles
-- Clock period (ns): 2
-- Target frequency (MHz): 500
-- Input signals: X Y Cin
-- Output signals: R
--  approx. input signal timings: X: (c0, 0.550000ns)Y: (c1, 1.110000ns)Cin: (c0, 0.000000ns)
--  approx. output signal timings: R: (c2, 0.610000ns)

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntAdder_30_Freq500_uid34 is
    port (clk : in std_logic;
          X : in  std_logic_vector(29 downto 0);
          Y : in  std_logic_vector(29 downto 0);
          Cin : in  std_logic;
          R : out  std_logic_vector(29 downto 0)   );
end entity;

architecture arch of IntAdder_30_Freq500_uid34 is
signal Cin_1, Cin_1_d1, Cin_1_d2 :  std_logic;
   -- timing of Cin_1: (c0, 0.000000ns)
signal X_1, X_1_d1, X_1_d2 :  std_logic_vector(30 downto 0);
   -- timing of X_1: (c0, 0.550000ns)
signal Y_1, Y_1_d1 :  std_logic_vector(30 downto 0);
   -- timing of Y_1: (c1, 1.110000ns)
signal S_1 :  std_logic_vector(30 downto 0);
   -- timing of S_1: (c2, 0.610000ns)
signal R_1 :  std_logic_vector(29 downto 0);
   -- timing of R_1: (c2, 0.610000ns)
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            Cin_1_d1 <=  Cin_1;
            Cin_1_d2 <=  Cin_1_d1;
            X_1_d1 <=  X_1;
            X_1_d2 <=  X_1_d1;
            Y_1_d1 <=  Y_1;
         end if;
      end process;
   Cin_1 <= Cin;
   X_1 <= '0' & X(29 downto 0);
   Y_1 <= '0' & Y(29 downto 0);
   S_1 <= X_1_d2 + Y_1_d1 + Cin_1_d2;
   R_1 <= S_1(29 downto 0);
   R <= R_1 ;
end architecture;

--------------------------------------------------------------------------------
--                         IntAdder_30_Freq500_uid37
-- VHDL generated for DummyFPGA @ 500MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin (2008-2016)
--------------------------------------------------------------------------------
-- Pipeline depth: 6 cycles
-- Clock period (ns): 2
-- Target frequency (MHz): 500
-- Input signals: X Y Cin
-- Output signals: R
--  approx. input signal timings: X: (c2, 0.610000ns)Y: (c6, 0.044615ns)Cin: (c0, 0.000000ns)
--  approx. output signal timings: R: (c6, 1.334615ns)

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntAdder_30_Freq500_uid37 is
    port (clk : in std_logic;
          X : in  std_logic_vector(29 downto 0);
          Y : in  std_logic_vector(29 downto 0);
          Cin : in  std_logic;
          R : out  std_logic_vector(29 downto 0)   );
end entity;

architecture arch of IntAdder_30_Freq500_uid37 is
signal Rtmp :  std_logic_vector(29 downto 0);
   -- timing of Rtmp: (c6, 1.334615ns)
signal X_d1, X_d2, X_d3, X_d4 :  std_logic_vector(29 downto 0);
   -- timing of X: (c2, 0.610000ns)
signal Cin_d1, Cin_d2, Cin_d3, Cin_d4, Cin_d5, Cin_d6 :  std_logic;
   -- timing of Cin: (c0, 0.000000ns)
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            X_d1 <=  X;
            X_d2 <=  X_d1;
            X_d3 <=  X_d2;
            X_d4 <=  X_d3;
            Cin_d1 <=  Cin;
            Cin_d2 <=  Cin_d1;
            Cin_d3 <=  Cin_d2;
            Cin_d4 <=  Cin_d3;
            Cin_d5 <=  Cin_d4;
            Cin_d6 <=  Cin_d5;
         end if;
      end process;
   Rtmp <= X_d4 + Y + Cin_d6;
   R <= Rtmp;
end architecture;

--------------------------------------------------------------------------------
--                         IntAdder_29_Freq500_uid49
-- VHDL generated for DummyFPGA @ 500MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin (2008-2016)
--------------------------------------------------------------------------------
-- Pipeline depth: 1 cycles
-- Clock period (ns): 2
-- Target frequency (MHz): 500
-- Input signals: X Y Cin
-- Output signals: R
--  approx. input signal timings: X: (c1, 0.370000ns)Y: (c1, 0.370000ns)Cin: (c0, 0.000000ns)
--  approx. output signal timings: R: (c1, 1.650000ns)

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntAdder_29_Freq500_uid49 is
    port (clk : in std_logic;
          X : in  std_logic_vector(28 downto 0);
          Y : in  std_logic_vector(28 downto 0);
          Cin : in  std_logic;
          R : out  std_logic_vector(28 downto 0)   );
end entity;

architecture arch of IntAdder_29_Freq500_uid49 is
signal Rtmp :  std_logic_vector(28 downto 0);
   -- timing of Rtmp: (c1, 1.650000ns)
signal Cin_d1 :  std_logic;
   -- timing of Cin: (c0, 0.000000ns)
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            Cin_d1 <=  Cin;
         end if;
      end process;
   Rtmp <= X + Y + Cin_d1;
   R <= Rtmp;
end architecture;

--------------------------------------------------------------------------------
--                          FixRealKCM_Freq500_uid39
-- VHDL generated for DummyFPGA @ 500MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin (2007-2016)
--------------------------------------------------------------------------------
-- Pipeline depth: 1 cycles
-- Clock period (ns): 2
-- Target frequency (MHz): 500
-- Input signals: X
-- Output signals: R
--  approx. input signal timings: X: (c0, 1.620000ns)
--  approx. output signal timings: R: (c1, 1.650000ns)

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity FixRealKCM_Freq500_uid39 is
    port (clk : in std_logic;
          X : in  std_logic_vector(7 downto 0);
          R : out  std_logic_vector(28 downto 0)   );
end entity;

architecture arch of FixRealKCM_Freq500_uid39 is
   component FixRealKCM_Freq500_uid39_T0_Freq500_uid42 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(28 downto 0)   );
   end component;

   component FixRealKCM_Freq500_uid39_T1_Freq500_uid45 is
      port ( X : in  std_logic_vector(2 downto 0);
             Y : out  std_logic_vector(23 downto 0)   );
   end component;

   component IntAdder_29_Freq500_uid49 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(28 downto 0);
             Y : in  std_logic_vector(28 downto 0);
             Cin : in  std_logic;
             R : out  std_logic_vector(28 downto 0)   );
   end component;

signal FixRealKCM_Freq500_uid39_A0 :  std_logic_vector(4 downto 0);
   -- timing of FixRealKCM_Freq500_uid39_A0: (c0, 1.620000ns)
signal FixRealKCM_Freq500_uid39_T0 :  std_logic_vector(28 downto 0);
   -- timing of FixRealKCM_Freq500_uid39_T0: (c1, 0.370000ns)
signal FixRealKCM_Freq500_uid39_T0_copy43, FixRealKCM_Freq500_uid39_T0_copy43_d1 :  std_logic_vector(28 downto 0);
   -- timing of FixRealKCM_Freq500_uid39_T0_copy43: (c0, 1.620000ns)
signal bh40_w0_0 :  std_logic;
   -- timing of bh40_w0_0: (c1, 0.370000ns)
signal bh40_w1_0 :  std_logic;
   -- timing of bh40_w1_0: (c1, 0.370000ns)
signal bh40_w2_0 :  std_logic;
   -- timing of bh40_w2_0: (c1, 0.370000ns)
signal bh40_w3_0 :  std_logic;
   -- timing of bh40_w3_0: (c1, 0.370000ns)
signal bh40_w4_0 :  std_logic;
   -- timing of bh40_w4_0: (c1, 0.370000ns)
signal bh40_w5_0 :  std_logic;
   -- timing of bh40_w5_0: (c1, 0.370000ns)
signal bh40_w6_0 :  std_logic;
   -- timing of bh40_w6_0: (c1, 0.370000ns)
signal bh40_w7_0 :  std_logic;
   -- timing of bh40_w7_0: (c1, 0.370000ns)
signal bh40_w8_0 :  std_logic;
   -- timing of bh40_w8_0: (c1, 0.370000ns)
signal bh40_w9_0 :  std_logic;
   -- timing of bh40_w9_0: (c1, 0.370000ns)
signal bh40_w10_0 :  std_logic;
   -- timing of bh40_w10_0: (c1, 0.370000ns)
signal bh40_w11_0 :  std_logic;
   -- timing of bh40_w11_0: (c1, 0.370000ns)
signal bh40_w12_0 :  std_logic;
   -- timing of bh40_w12_0: (c1, 0.370000ns)
signal bh40_w13_0 :  std_logic;
   -- timing of bh40_w13_0: (c1, 0.370000ns)
signal bh40_w14_0 :  std_logic;
   -- timing of bh40_w14_0: (c1, 0.370000ns)
signal bh40_w15_0 :  std_logic;
   -- timing of bh40_w15_0: (c1, 0.370000ns)
signal bh40_w16_0 :  std_logic;
   -- timing of bh40_w16_0: (c1, 0.370000ns)
signal bh40_w17_0 :  std_logic;
   -- timing of bh40_w17_0: (c1, 0.370000ns)
signal bh40_w18_0 :  std_logic;
   -- timing of bh40_w18_0: (c1, 0.370000ns)
signal bh40_w19_0 :  std_logic;
   -- timing of bh40_w19_0: (c1, 0.370000ns)
signal bh40_w20_0 :  std_logic;
   -- timing of bh40_w20_0: (c1, 0.370000ns)
signal bh40_w21_0 :  std_logic;
   -- timing of bh40_w21_0: (c1, 0.370000ns)
signal bh40_w22_0 :  std_logic;
   -- timing of bh40_w22_0: (c1, 0.370000ns)
signal bh40_w23_0 :  std_logic;
   -- timing of bh40_w23_0: (c1, 0.370000ns)
signal bh40_w24_0 :  std_logic;
   -- timing of bh40_w24_0: (c1, 0.370000ns)
signal bh40_w25_0 :  std_logic;
   -- timing of bh40_w25_0: (c1, 0.370000ns)
signal bh40_w26_0 :  std_logic;
   -- timing of bh40_w26_0: (c1, 0.370000ns)
signal bh40_w27_0 :  std_logic;
   -- timing of bh40_w27_0: (c1, 0.370000ns)
signal bh40_w28_0 :  std_logic;
   -- timing of bh40_w28_0: (c1, 0.370000ns)
signal FixRealKCM_Freq500_uid39_A1 :  std_logic_vector(2 downto 0);
   -- timing of FixRealKCM_Freq500_uid39_A1: (c0, 1.620000ns)
signal FixRealKCM_Freq500_uid39_T1 :  std_logic_vector(23 downto 0);
   -- timing of FixRealKCM_Freq500_uid39_T1: (c1, 0.370000ns)
signal FixRealKCM_Freq500_uid39_T1_copy46, FixRealKCM_Freq500_uid39_T1_copy46_d1 :  std_logic_vector(23 downto 0);
   -- timing of FixRealKCM_Freq500_uid39_T1_copy46: (c0, 1.620000ns)
signal bh40_w0_1 :  std_logic;
   -- timing of bh40_w0_1: (c1, 0.370000ns)
signal bh40_w1_1 :  std_logic;
   -- timing of bh40_w1_1: (c1, 0.370000ns)
signal bh40_w2_1 :  std_logic;
   -- timing of bh40_w2_1: (c1, 0.370000ns)
signal bh40_w3_1 :  std_logic;
   -- timing of bh40_w3_1: (c1, 0.370000ns)
signal bh40_w4_1 :  std_logic;
   -- timing of bh40_w4_1: (c1, 0.370000ns)
signal bh40_w5_1 :  std_logic;
   -- timing of bh40_w5_1: (c1, 0.370000ns)
signal bh40_w6_1 :  std_logic;
   -- timing of bh40_w6_1: (c1, 0.370000ns)
signal bh40_w7_1 :  std_logic;
   -- timing of bh40_w7_1: (c1, 0.370000ns)
signal bh40_w8_1 :  std_logic;
   -- timing of bh40_w8_1: (c1, 0.370000ns)
signal bh40_w9_1 :  std_logic;
   -- timing of bh40_w9_1: (c1, 0.370000ns)
signal bh40_w10_1 :  std_logic;
   -- timing of bh40_w10_1: (c1, 0.370000ns)
signal bh40_w11_1 :  std_logic;
   -- timing of bh40_w11_1: (c1, 0.370000ns)
signal bh40_w12_1 :  std_logic;
   -- timing of bh40_w12_1: (c1, 0.370000ns)
signal bh40_w13_1 :  std_logic;
   -- timing of bh40_w13_1: (c1, 0.370000ns)
signal bh40_w14_1 :  std_logic;
   -- timing of bh40_w14_1: (c1, 0.370000ns)
signal bh40_w15_1 :  std_logic;
   -- timing of bh40_w15_1: (c1, 0.370000ns)
signal bh40_w16_1 :  std_logic;
   -- timing of bh40_w16_1: (c1, 0.370000ns)
signal bh40_w17_1 :  std_logic;
   -- timing of bh40_w17_1: (c1, 0.370000ns)
signal bh40_w18_1 :  std_logic;
   -- timing of bh40_w18_1: (c1, 0.370000ns)
signal bh40_w19_1 :  std_logic;
   -- timing of bh40_w19_1: (c1, 0.370000ns)
signal bh40_w20_1 :  std_logic;
   -- timing of bh40_w20_1: (c1, 0.370000ns)
signal bh40_w21_1 :  std_logic;
   -- timing of bh40_w21_1: (c1, 0.370000ns)
signal bh40_w22_1 :  std_logic;
   -- timing of bh40_w22_1: (c1, 0.370000ns)
signal bh40_w23_1 :  std_logic;
   -- timing of bh40_w23_1: (c1, 0.370000ns)
signal bitheapFinalAdd_bh40_In0 :  std_logic_vector(28 downto 0);
   -- timing of bitheapFinalAdd_bh40_In0: (c1, 0.370000ns)
signal bitheapFinalAdd_bh40_In1 :  std_logic_vector(28 downto 0);
   -- timing of bitheapFinalAdd_bh40_In1: (c1, 0.370000ns)
signal bitheapFinalAdd_bh40_Cin :  std_logic;
   -- timing of bitheapFinalAdd_bh40_Cin: (c0, 0.000000ns)
signal bitheapFinalAdd_bh40_Out :  std_logic_vector(28 downto 0);
   -- timing of bitheapFinalAdd_bh40_Out: (c1, 1.650000ns)
signal bitheapResult_bh40 :  std_logic_vector(28 downto 0);
   -- timing of bitheapResult_bh40: (c1, 1.650000ns)
signal OutRes :  std_logic_vector(28 downto 0);
   -- timing of OutRes: (c1, 1.650000ns)
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            FixRealKCM_Freq500_uid39_T0_copy43_d1 <=  FixRealKCM_Freq500_uid39_T0_copy43;
            FixRealKCM_Freq500_uid39_T1_copy46_d1 <=  FixRealKCM_Freq500_uid39_T1_copy46;
         end if;
      end process;
-- This operator multiplies by log(2)
   FixRealKCM_Freq500_uid39_A0 <= X(7 downto 3);-- input address  m=7  l=3
   FixRealKCM_Freq500_uid39_Table0: FixRealKCM_Freq500_uid39_T0_Freq500_uid42
      port map ( X => FixRealKCM_Freq500_uid39_A0,
                 Y => FixRealKCM_Freq500_uid39_T0_copy43);
   FixRealKCM_Freq500_uid39_T0 <= FixRealKCM_Freq500_uid39_T0_copy43_d1; -- output copy to hold a pipeline register if needed
   bh40_w0_0 <= FixRealKCM_Freq500_uid39_T0(0);
   bh40_w1_0 <= FixRealKCM_Freq500_uid39_T0(1);
   bh40_w2_0 <= FixRealKCM_Freq500_uid39_T0(2);
   bh40_w3_0 <= FixRealKCM_Freq500_uid39_T0(3);
   bh40_w4_0 <= FixRealKCM_Freq500_uid39_T0(4);
   bh40_w5_0 <= FixRealKCM_Freq500_uid39_T0(5);
   bh40_w6_0 <= FixRealKCM_Freq500_uid39_T0(6);
   bh40_w7_0 <= FixRealKCM_Freq500_uid39_T0(7);
   bh40_w8_0 <= FixRealKCM_Freq500_uid39_T0(8);
   bh40_w9_0 <= FixRealKCM_Freq500_uid39_T0(9);
   bh40_w10_0 <= FixRealKCM_Freq500_uid39_T0(10);
   bh40_w11_0 <= FixRealKCM_Freq500_uid39_T0(11);
   bh40_w12_0 <= FixRealKCM_Freq500_uid39_T0(12);
   bh40_w13_0 <= FixRealKCM_Freq500_uid39_T0(13);
   bh40_w14_0 <= FixRealKCM_Freq500_uid39_T0(14);
   bh40_w15_0 <= FixRealKCM_Freq500_uid39_T0(15);
   bh40_w16_0 <= FixRealKCM_Freq500_uid39_T0(16);
   bh40_w17_0 <= FixRealKCM_Freq500_uid39_T0(17);
   bh40_w18_0 <= FixRealKCM_Freq500_uid39_T0(18);
   bh40_w19_0 <= FixRealKCM_Freq500_uid39_T0(19);
   bh40_w20_0 <= FixRealKCM_Freq500_uid39_T0(20);
   bh40_w21_0 <= FixRealKCM_Freq500_uid39_T0(21);
   bh40_w22_0 <= FixRealKCM_Freq500_uid39_T0(22);
   bh40_w23_0 <= FixRealKCM_Freq500_uid39_T0(23);
   bh40_w24_0 <= FixRealKCM_Freq500_uid39_T0(24);
   bh40_w25_0 <= FixRealKCM_Freq500_uid39_T0(25);
   bh40_w26_0 <= FixRealKCM_Freq500_uid39_T0(26);
   bh40_w27_0 <= FixRealKCM_Freq500_uid39_T0(27);
   bh40_w28_0 <= FixRealKCM_Freq500_uid39_T0(28);
   FixRealKCM_Freq500_uid39_A1 <= X(2 downto 0);-- input address  m=2  l=0
   FixRealKCM_Freq500_uid39_Table1: FixRealKCM_Freq500_uid39_T1_Freq500_uid45
      port map ( X => FixRealKCM_Freq500_uid39_A1,
                 Y => FixRealKCM_Freq500_uid39_T1_copy46);
   FixRealKCM_Freq500_uid39_T1 <= FixRealKCM_Freq500_uid39_T1_copy46_d1; -- output copy to hold a pipeline register if needed
   bh40_w0_1 <= FixRealKCM_Freq500_uid39_T1(0);
   bh40_w1_1 <= FixRealKCM_Freq500_uid39_T1(1);
   bh40_w2_1 <= FixRealKCM_Freq500_uid39_T1(2);
   bh40_w3_1 <= FixRealKCM_Freq500_uid39_T1(3);
   bh40_w4_1 <= FixRealKCM_Freq500_uid39_T1(4);
   bh40_w5_1 <= FixRealKCM_Freq500_uid39_T1(5);
   bh40_w6_1 <= FixRealKCM_Freq500_uid39_T1(6);
   bh40_w7_1 <= FixRealKCM_Freq500_uid39_T1(7);
   bh40_w8_1 <= FixRealKCM_Freq500_uid39_T1(8);
   bh40_w9_1 <= FixRealKCM_Freq500_uid39_T1(9);
   bh40_w10_1 <= FixRealKCM_Freq500_uid39_T1(10);
   bh40_w11_1 <= FixRealKCM_Freq500_uid39_T1(11);
   bh40_w12_1 <= FixRealKCM_Freq500_uid39_T1(12);
   bh40_w13_1 <= FixRealKCM_Freq500_uid39_T1(13);
   bh40_w14_1 <= FixRealKCM_Freq500_uid39_T1(14);
   bh40_w15_1 <= FixRealKCM_Freq500_uid39_T1(15);
   bh40_w16_1 <= FixRealKCM_Freq500_uid39_T1(16);
   bh40_w17_1 <= FixRealKCM_Freq500_uid39_T1(17);
   bh40_w18_1 <= FixRealKCM_Freq500_uid39_T1(18);
   bh40_w19_1 <= FixRealKCM_Freq500_uid39_T1(19);
   bh40_w20_1 <= FixRealKCM_Freq500_uid39_T1(20);
   bh40_w21_1 <= FixRealKCM_Freq500_uid39_T1(21);
   bh40_w22_1 <= FixRealKCM_Freq500_uid39_T1(22);
   bh40_w23_1 <= FixRealKCM_Freq500_uid39_T1(23);

   -- Adding the constant bits 
      -- All the constant bits are zero, nothing to add


   bitheapFinalAdd_bh40_In0 <= "" & bh40_w28_0 & bh40_w27_0 & bh40_w26_0 & bh40_w25_0 & bh40_w24_0 & bh40_w23_1 & bh40_w22_1 & bh40_w21_1 & bh40_w20_1 & bh40_w19_1 & bh40_w18_1 & bh40_w17_1 & bh40_w16_1 & bh40_w15_1 & bh40_w14_1 & bh40_w13_1 & bh40_w12_1 & bh40_w11_1 & bh40_w10_1 & bh40_w9_1 & bh40_w8_1 & bh40_w7_1 & bh40_w6_1 & bh40_w5_1 & bh40_w4_1 & bh40_w3_1 & bh40_w2_1 & bh40_w1_1 & bh40_w0_1;
   bitheapFinalAdd_bh40_In1 <= "0" & "0" & "0" & "0" & "0" & bh40_w23_0 & bh40_w22_0 & bh40_w21_0 & bh40_w20_0 & bh40_w19_0 & bh40_w18_0 & bh40_w17_0 & bh40_w16_0 & bh40_w15_0 & bh40_w14_0 & bh40_w13_0 & bh40_w12_0 & bh40_w11_0 & bh40_w10_0 & bh40_w9_0 & bh40_w8_0 & bh40_w7_0 & bh40_w6_0 & bh40_w5_0 & bh40_w4_0 & bh40_w3_0 & bh40_w2_0 & bh40_w1_0 & bh40_w0_0;
   bitheapFinalAdd_bh40_Cin <= '0';

   bitheapFinalAdd_bh40: IntAdder_29_Freq500_uid49
      port map ( clk  => clk,
                 Cin => bitheapFinalAdd_bh40_Cin,
                 X => bitheapFinalAdd_bh40_In0,
                 Y => bitheapFinalAdd_bh40_In1,
                 R => bitheapFinalAdd_bh40_Out);
   bitheapResult_bh40 <= bitheapFinalAdd_bh40_Out(28 downto 0);
   OutRes <= bitheapResult_bh40(28 downto 0);
   R <= OutRes(28 downto 0);
end architecture;

--------------------------------------------------------------------------------
--                         IntAdder_38_Freq500_uid51
-- VHDL generated for DummyFPGA @ 500MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin (2008-2016)
--------------------------------------------------------------------------------
-- Pipeline depth: 8 cycles
-- Clock period (ns): 2
-- Target frequency (MHz): 500
-- Input signals: X Y Cin
-- Output signals: R
--  approx. input signal timings: X: (c1, 1.650000ns)Y: (c6, 1.334615ns)Cin: (c0, 0.550000ns)
--  approx. output signal timings: R: (c8, 0.114615ns)

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntAdder_38_Freq500_uid51 is
    port (clk : in std_logic;
          X : in  std_logic_vector(37 downto 0);
          Y : in  std_logic_vector(37 downto 0);
          Cin : in  std_logic;
          R : out  std_logic_vector(37 downto 0)   );
end entity;

architecture arch of IntAdder_38_Freq500_uid51 is
signal Cin_0, Cin_0_d1, Cin_0_d2, Cin_0_d3, Cin_0_d4, Cin_0_d5, Cin_0_d6, Cin_0_d7 :  std_logic;
   -- timing of Cin_0: (c0, 0.550000ns)
signal X_0, X_0_d1, X_0_d2, X_0_d3, X_0_d4, X_0_d5, X_0_d6 :  std_logic_vector(25 downto 0);
   -- timing of X_0: (c1, 1.650000ns)
signal Y_0, Y_0_d1 :  std_logic_vector(25 downto 0);
   -- timing of Y_0: (c6, 1.334615ns)
signal S_0 :  std_logic_vector(25 downto 0);
   -- timing of S_0: (c7, 0.784615ns)
signal R_0, R_0_d1 :  std_logic_vector(24 downto 0);
   -- timing of R_0: (c7, 0.784615ns)
signal Cin_1, Cin_1_d1 :  std_logic;
   -- timing of Cin_1: (c7, 0.784615ns)
signal X_1, X_1_d1, X_1_d2, X_1_d3, X_1_d4, X_1_d5, X_1_d6, X_1_d7 :  std_logic_vector(13 downto 0);
   -- timing of X_1: (c1, 1.650000ns)
signal Y_1, Y_1_d1, Y_1_d2 :  std_logic_vector(13 downto 0);
   -- timing of Y_1: (c6, 1.334615ns)
signal S_1 :  std_logic_vector(13 downto 0);
   -- timing of S_1: (c8, 0.114615ns)
signal R_1 :  std_logic_vector(12 downto 0);
   -- timing of R_1: (c8, 0.114615ns)
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            Cin_0_d1 <=  Cin_0;
            Cin_0_d2 <=  Cin_0_d1;
            Cin_0_d3 <=  Cin_0_d2;
            Cin_0_d4 <=  Cin_0_d3;
            Cin_0_d5 <=  Cin_0_d4;
            Cin_0_d6 <=  Cin_0_d5;
            Cin_0_d7 <=  Cin_0_d6;
            X_0_d1 <=  X_0;
            X_0_d2 <=  X_0_d1;
            X_0_d3 <=  X_0_d2;
            X_0_d4 <=  X_0_d3;
            X_0_d5 <=  X_0_d4;
            X_0_d6 <=  X_0_d5;
            Y_0_d1 <=  Y_0;
            R_0_d1 <=  R_0;
            Cin_1_d1 <=  Cin_1;
            X_1_d1 <=  X_1;
            X_1_d2 <=  X_1_d1;
            X_1_d3 <=  X_1_d2;
            X_1_d4 <=  X_1_d3;
            X_1_d5 <=  X_1_d4;
            X_1_d6 <=  X_1_d5;
            X_1_d7 <=  X_1_d6;
            Y_1_d1 <=  Y_1;
            Y_1_d2 <=  Y_1_d1;
         end if;
      end process;
   Cin_0 <= Cin;
   X_0 <= '0' & X(24 downto 0);
   Y_0 <= '0' & Y(24 downto 0);
   S_0 <= X_0_d6 + Y_0_d1 + Cin_0_d7;
   R_0 <= S_0(24 downto 0);
   Cin_1 <= S_0(25);
   X_1 <= '0' & X(37 downto 25);
   Y_1 <= '0' & Y(37 downto 25);
   S_1 <= X_1_d7 + Y_1_d2 + Cin_1_d1;
   R_1 <= S_1(12 downto 0);
   R <= R_1 & R_0_d1 ;
end architecture;

--------------------------------------------------------------------------------
--                    Normalizer_Z_38_30_16_Freq500_uid53
-- VHDL generated for DummyFPGA @ 500MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, (2007-2020)
--------------------------------------------------------------------------------
-- Pipeline depth: 3 cycles
-- Clock period (ns): 2
-- Target frequency (MHz): 500
-- Input signals: X
-- Output signals: Count R
--  approx. input signal timings: X: (c8, 0.114615ns)
--  approx. output signal timings: Count: (c10, 1.554615ns)R: (c11, 0.304615ns)

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity Normalizer_Z_38_30_16_Freq500_uid53 is
    port (clk : in std_logic;
          X : in  std_logic_vector(37 downto 0);
          Count : out  std_logic_vector(4 downto 0);
          R : out  std_logic_vector(29 downto 0)   );
end entity;

architecture arch of Normalizer_Z_38_30_16_Freq500_uid53 is
signal level5 :  std_logic_vector(37 downto 0);
   -- timing of level5: (c8, 0.114615ns)
signal count4, count4_d1, count4_d2 :  std_logic;
   -- timing of count4: (c8, 0.704615ns)
signal level4, level4_d1 :  std_logic_vector(37 downto 0);
   -- timing of level4: (c8, 1.254615ns)
signal count3, count3_d1 :  std_logic;
   -- timing of count3: (c9, 0.024615ns)
signal level3 :  std_logic_vector(36 downto 0);
   -- timing of level3: (c9, 0.574615ns)
signal count2, count2_d1 :  std_logic;
   -- timing of count2: (c9, 1.134615ns)
signal level2, level2_d1 :  std_logic_vector(32 downto 0);
   -- timing of level2: (c9, 1.684615ns)
signal count1 :  std_logic;
   -- timing of count1: (c10, 0.444615ns)
signal level1, level1_d1 :  std_logic_vector(30 downto 0);
   -- timing of level1: (c10, 0.994615ns)
signal count0, count0_d1 :  std_logic;
   -- timing of count0: (c10, 1.554615ns)
signal level0 :  std_logic_vector(29 downto 0);
   -- timing of level0: (c11, 0.304615ns)
signal sCount :  std_logic_vector(4 downto 0);
   -- timing of sCount: (c10, 1.554615ns)
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            count4_d1 <=  count4;
            count4_d2 <=  count4_d1;
            level4_d1 <=  level4;
            count3_d1 <=  count3;
            count2_d1 <=  count2;
            level2_d1 <=  level2;
            level1_d1 <=  level1;
            count0_d1 <=  count0;
         end if;
      end process;
   level5 <= X ;
   count4<= '1' when level5(37 downto 22) = (37 downto 22=>'0') else '0';
   level4<= level5(37 downto 0) when count4='0' else level5(21 downto 0) & (15 downto 0 => '0');

   count3<= '1' when level4_d1(37 downto 30) = (37 downto 30=>'0') else '0';
   level3<= level4_d1(37 downto 1) when count3='0' else level4_d1(29 downto 0) & (6 downto 0 => '0');

   count2<= '1' when level3(36 downto 33) = (36 downto 33=>'0') else '0';
   level2<= level3(36 downto 4) when count2='0' else level3(32 downto 0);

   count1<= '1' when level2_d1(32 downto 31) = (32 downto 31=>'0') else '0';
   level1<= level2_d1(32 downto 2) when count1='0' else level2_d1(30 downto 0);

   count0<= '1' when level1(30 downto 30) = (30 downto 30=>'0') else '0';
   level0<= level1_d1(30 downto 1) when count0_d1='0' else level1_d1(29 downto 0);

   R <= level0;
   sCount <= count4_d2 & count3_d1 & count2_d1 & count1 & count0;
   Count <= sCount;
end architecture;

--------------------------------------------------------------------------------
--                   RightShifter14_by_max_13_Freq500_uid55
-- VHDL generated for DummyFPGA @ 500MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca (2008-2011), Florent de Dinechin (2008-2019)
--------------------------------------------------------------------------------
-- Pipeline depth: 3 cycles
-- Clock period (ns): 2
-- Target frequency (MHz): 500
-- Input signals: X S
-- Output signals: R
--  approx. input signal timings: X: (c5, 0.094615ns)S: (c3, 1.460000ns)
--  approx. output signal timings: R: (c6, 0.102308ns)

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity RightShifter14_by_max_13_Freq500_uid55 is
    port (clk : in std_logic;
          X : in  std_logic_vector(13 downto 0);
          S : in  std_logic_vector(3 downto 0);
          R : out  std_logic_vector(26 downto 0)   );
end entity;

architecture arch of RightShifter14_by_max_13_Freq500_uid55 is
signal ps, ps_d1, ps_d2, ps_d3 :  std_logic_vector(3 downto 0);
   -- timing of ps: (c3, 1.460000ns)
signal level0 :  std_logic_vector(13 downto 0);
   -- timing of level0: (c5, 0.094615ns)
signal level1 :  std_logic_vector(14 downto 0);
   -- timing of level1: (c5, 0.094615ns)
signal level2 :  std_logic_vector(16 downto 0);
   -- timing of level2: (c5, 0.906154ns)
signal level3, level3_d1 :  std_logic_vector(20 downto 0);
   -- timing of level3: (c5, 0.906154ns)
signal level4 :  std_logic_vector(28 downto 0);
   -- timing of level4: (c6, 0.102308ns)
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            ps_d1 <=  ps;
            ps_d2 <=  ps_d1;
            ps_d3 <=  ps_d2;
            level3_d1 <=  level3;
         end if;
      end process;
   ps<= S;
   level0<= X;
   level1 <=  (0 downto 0 => '0') & level0 when ps_d2(0) = '1' else    level0 & (0 downto 0 => '0');
   level2 <=  (1 downto 0 => '0') & level1 when ps_d2(1) = '1' else    level1 & (1 downto 0 => '0');
   level3 <=  (3 downto 0 => '0') & level2 when ps_d2(2) = '1' else    level2 & (3 downto 0 => '0');
   level4 <=  (7 downto 0 => '0') & level3_d1 when ps_d3(3) = '1' else    level3_d1 & (7 downto 0 => '0');
   R <= level4(28 downto 2);
end architecture;

--------------------------------------------------------------------------------
--                         IntAdder_23_Freq500_uid57
-- VHDL generated for DummyFPGA @ 500MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin (2008-2016)
--------------------------------------------------------------------------------
-- Pipeline depth: 6 cycles
-- Clock period (ns): 2
-- Target frequency (MHz): 500
-- Input signals: X Y Cin
-- Output signals: R
--  approx. input signal timings: X: (c4, 1.344615ns)Y: (c6, 0.102308ns)Cin: (c0, 0.550000ns)
--  approx. output signal timings: R: (c6, 1.322308ns)

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntAdder_23_Freq500_uid57 is
    port (clk : in std_logic;
          X : in  std_logic_vector(22 downto 0);
          Y : in  std_logic_vector(22 downto 0);
          Cin : in  std_logic;
          R : out  std_logic_vector(22 downto 0)   );
end entity;

architecture arch of IntAdder_23_Freq500_uid57 is
signal Rtmp :  std_logic_vector(22 downto 0);
   -- timing of Rtmp: (c6, 1.322308ns)
signal X_d1, X_d2 :  std_logic_vector(22 downto 0);
   -- timing of X: (c4, 1.344615ns)
signal Cin_d1, Cin_d2, Cin_d3, Cin_d4, Cin_d5, Cin_d6 :  std_logic;
   -- timing of Cin: (c0, 0.550000ns)
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            X_d1 <=  X;
            X_d2 <=  X_d1;
            Cin_d1 <=  Cin;
            Cin_d2 <=  Cin_d1;
            Cin_d3 <=  Cin_d2;
            Cin_d4 <=  Cin_d3;
            Cin_d5 <=  Cin_d4;
            Cin_d6 <=  Cin_d5;
         end if;
      end process;
   Rtmp <= X_d2 + Y + Cin_d6;
   R <= Rtmp;
end architecture;

--------------------------------------------------------------------------------
--                         IntAdder_25_Freq500_uid60
-- VHDL generated for DummyFPGA @ 500MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin (2008-2016)
--------------------------------------------------------------------------------
-- Pipeline depth: 11 cycles
-- Clock period (ns): 2
-- Target frequency (MHz): 500
-- Input signals: X Y Cin
-- Output signals: R
--  approx. input signal timings: X: (c11, 0.304615ns)Y: (c11, 0.304615ns)Cin: (c0, 0.000000ns)
--  approx. output signal timings: R: (c11, 1.544615ns)

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntAdder_25_Freq500_uid60 is
    port (clk : in std_logic;
          X : in  std_logic_vector(24 downto 0);
          Y : in  std_logic_vector(24 downto 0);
          Cin : in  std_logic;
          R : out  std_logic_vector(24 downto 0)   );
end entity;

architecture arch of IntAdder_25_Freq500_uid60 is
signal Rtmp :  std_logic_vector(24 downto 0);
   -- timing of Rtmp: (c11, 1.544615ns)
signal Cin_d1, Cin_d2, Cin_d3, Cin_d4, Cin_d5, Cin_d6, Cin_d7, Cin_d8, Cin_d9, Cin_d10, Cin_d11 :  std_logic;
   -- timing of Cin: (c0, 0.000000ns)
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            Cin_d1 <=  Cin;
            Cin_d2 <=  Cin_d1;
            Cin_d3 <=  Cin_d2;
            Cin_d4 <=  Cin_d3;
            Cin_d5 <=  Cin_d4;
            Cin_d6 <=  Cin_d5;
            Cin_d7 <=  Cin_d6;
            Cin_d8 <=  Cin_d7;
            Cin_d9 <=  Cin_d8;
            Cin_d10 <=  Cin_d9;
            Cin_d11 <=  Cin_d10;
         end if;
      end process;
   Rtmp <= X + Y + Cin_d11;
   R <= Rtmp;
end architecture;

--------------------------------------------------------------------------------
--                   FPLogIterative_8_17_0_500_Freq500_uid9
-- VHDL generated for DummyFPGA @ 500MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: F. de Dinechin, C. Klein  (2008-2011)
--------------------------------------------------------------------------------
-- Pipeline depth: 11 cycles
-- Clock period (ns): 2
-- Target frequency (MHz): 500
-- Input signals: X
-- Output signals: R
--  approx. input signal timings: X: (c0, 0.000000ns)
--  approx. output signal timings: R: (c11, 1.544615ns)

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity FPLogIterative_8_17_0_500_Freq500_uid9 is
    port (clk : in std_logic;
          X : in  std_logic_vector(8+17+2 downto 0);
          R : out  std_logic_vector(8+17+2 downto 0)   );
end entity;

architecture arch of FPLogIterative_8_17_0_500_Freq500_uid9 is
   component LZOC_17_Freq500_uid11 is
      port ( clk : in std_logic;
             I : in  std_logic_vector(16 downto 0);
             OZB : in  std_logic;
             O : out  std_logic_vector(4 downto 0)   );
   end component;

   component LeftShifter10_by_max_10_Freq500_uid13 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(9 downto 0);
             S : in  std_logic_vector(3 downto 0);
             R : out  std_logic_vector(19 downto 0)   );
   end component;

   component InvA0Table_Freq500_uid15 is
      port ( X : in  std_logic_vector(6 downto 0);
             Y : out  std_logic_vector(7 downto 0)   );
   end component;

   component IntAdder_21_Freq500_uid19 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(20 downto 0);
             Y : in  std_logic_vector(20 downto 0);
             Cin : in  std_logic;
             R : out  std_logic_vector(20 downto 0)   );
   end component;

   component IntAdder_21_Freq500_uid22 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(20 downto 0);
             Y : in  std_logic_vector(20 downto 0);
             Cin : in  std_logic;
             R : out  std_logic_vector(20 downto 0)   );
   end component;

   component IntAdder_21_Freq500_uid25 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(20 downto 0);
             Y : in  std_logic_vector(20 downto 0);
             Cin : in  std_logic;
             R : out  std_logic_vector(20 downto 0)   );
   end component;

   component LogTable0_Freq500_uid27 is
      port ( X : in  std_logic_vector(6 downto 0);
             Y : out  std_logic_vector(29 downto 0)   );
   end component;

   component LogTable1_Freq500_uid30 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(24 downto 0)   );
   end component;

   component IntAdder_30_Freq500_uid34 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(29 downto 0);
             Y : in  std_logic_vector(29 downto 0);
             Cin : in  std_logic;
             R : out  std_logic_vector(29 downto 0)   );
   end component;

   component IntAdder_30_Freq500_uid37 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(29 downto 0);
             Y : in  std_logic_vector(29 downto 0);
             Cin : in  std_logic;
             R : out  std_logic_vector(29 downto 0)   );
   end component;

   component FixRealKCM_Freq500_uid39 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(7 downto 0);
             R : out  std_logic_vector(28 downto 0)   );
   end component;

   component IntAdder_38_Freq500_uid51 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(37 downto 0);
             Y : in  std_logic_vector(37 downto 0);
             Cin : in  std_logic;
             R : out  std_logic_vector(37 downto 0)   );
   end component;

   component Normalizer_Z_38_30_16_Freq500_uid53 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(37 downto 0);
             Count : out  std_logic_vector(4 downto 0);
             R : out  std_logic_vector(29 downto 0)   );
   end component;

   component RightShifter14_by_max_13_Freq500_uid55 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(13 downto 0);
             S : in  std_logic_vector(3 downto 0);
             R : out  std_logic_vector(26 downto 0)   );
   end component;

   component IntAdder_23_Freq500_uid57 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(22 downto 0);
             Y : in  std_logic_vector(22 downto 0);
             Cin : in  std_logic;
             R : out  std_logic_vector(22 downto 0)   );
   end component;

   component IntAdder_25_Freq500_uid60 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(24 downto 0);
             Y : in  std_logic_vector(24 downto 0);
             Cin : in  std_logic;
             R : out  std_logic_vector(24 downto 0)   );
   end component;

signal XExnSgn, XExnSgn_d1, XExnSgn_d2, XExnSgn_d3, XExnSgn_d4, XExnSgn_d5, XExnSgn_d6, XExnSgn_d7, XExnSgn_d8, XExnSgn_d9, XExnSgn_d10, XExnSgn_d11 :  std_logic_vector(2 downto 0);
   -- timing of XExnSgn: (c0, 0.000000ns)
signal FirstBit :  std_logic;
   -- timing of FirstBit: (c0, 0.000000ns)
signal Y0, Y0_d1 :  std_logic_vector(18 downto 0);
   -- timing of Y0: (c0, 0.550000ns)
signal Y0h :  std_logic_vector(16 downto 0);
   -- timing of Y0h: (c0, 0.550000ns)
signal sR, sR_d1, sR_d2, sR_d3, sR_d4, sR_d5, sR_d6, sR_d7, sR_d8, sR_d9, sR_d10, sR_d11 :  std_logic;
   -- timing of sR: (c0, 0.550000ns)
signal absZ0 :  std_logic_vector(9 downto 0);
   -- timing of absZ0: (c0, 1.640000ns)
signal E :  std_logic_vector(7 downto 0);
   -- timing of E: (c0, 1.070000ns)
signal absE :  std_logic_vector(7 downto 0);
   -- timing of absE: (c0, 1.620000ns)
signal EeqZero, EeqZero_d1, EeqZero_d2, EeqZero_d3, EeqZero_d4 :  std_logic;
   -- timing of EeqZero: (c0, 1.620000ns)
signal lzo, lzo_d1, lzo_d2, lzo_d3 :  std_logic_vector(4 downto 0);
   -- timing of lzo: (c3, 0.410000ns)
signal pfinal_s, pfinal_s_d1, pfinal_s_d2, pfinal_s_d3 :  std_logic_vector(4 downto 0);
   -- timing of pfinal_s: (c0, 0.000000ns)
signal shiftval :  std_logic_vector(5 downto 0);
   -- timing of shiftval: (c3, 1.460000ns)
signal shiftvalinL :  std_logic_vector(3 downto 0);
   -- timing of shiftvalinL: (c3, 1.460000ns)
signal shiftvalinR :  std_logic_vector(3 downto 0);
   -- timing of shiftvalinR: (c3, 1.460000ns)
signal doRR, doRR_d1, doRR_d2 :  std_logic;
   -- timing of doRR: (c3, 1.460000ns)
signal small, small_d1, small_d2, small_d3, small_d4, small_d5, small_d6, small_d7 :  std_logic;
   -- timing of small: (c4, 0.210000ns)
signal small_absZ0_normd_full :  std_logic_vector(19 downto 0);
   -- timing of small_absZ0_normd_full: (c4, 1.344615ns)
signal small_absZ0_normd, small_absZ0_normd_d1 :  std_logic_vector(9 downto 0);
   -- timing of small_absZ0_normd: (c4, 1.344615ns)
signal A0 :  std_logic_vector(6 downto 0);
   -- timing of A0: (c0, 0.000000ns)
signal InvA0, InvA0_d1 :  std_logic_vector(7 downto 0);
   -- timing of InvA0: (c0, 0.550000ns)
signal InvA0_copy16 :  std_logic_vector(7 downto 0);
   -- timing of InvA0_copy16: (c0, 0.000000ns)
signal P0 :  std_logic_vector(26 downto 0);
   -- timing of P0: (c1, 0.560000ns)
signal Z1 :  std_logic_vector(19 downto 0);
   -- timing of Z1: (c1, 0.560000ns)
signal A1, A1_d1 :  std_logic_vector(4 downto 0);
   -- timing of A1: (c1, 0.560000ns)
signal B1 :  std_logic_vector(14 downto 0);
   -- timing of B1: (c1, 0.560000ns)
signal ZM1, ZM1_d1 :  std_logic_vector(19 downto 0);
   -- timing of ZM1: (c1, 0.560000ns)
signal P1 :  std_logic_vector(24 downto 0);
   -- timing of P1: (c2, 0.550000ns)
signal Y1 :  std_logic_vector(25 downto 0);
   -- timing of Y1: (c1, 0.560000ns)
signal EiY1 :  std_logic_vector(20 downto 0);
   -- timing of EiY1: (c1, 1.110000ns)
signal addXIter1 :  std_logic_vector(20 downto 0);
   -- timing of addXIter1: (c1, 0.560000ns)
signal EiYPB1 :  std_logic_vector(20 downto 0);
   -- timing of EiYPB1: (c2, 0.520000ns)
signal Pp1 :  std_logic_vector(20 downto 0);
   -- timing of Pp1: (c2, 1.100000ns)
signal Z2 :  std_logic_vector(20 downto 0);
   -- timing of Z2: (c3, 0.510000ns)
signal Zfinal, Zfinal_d1, Zfinal_d2 :  std_logic_vector(20 downto 0);
   -- timing of Zfinal: (c3, 0.510000ns)
signal squarerIn :  std_logic_vector(13 downto 0);
   -- timing of squarerIn: (c5, 0.094615ns)
signal Z2o2_full :  std_logic_vector(27 downto 0);
   -- timing of Z2o2_full: (c5, 0.094615ns)
signal Z2o2_full_dummy :  std_logic_vector(27 downto 0);
   -- timing of Z2o2_full_dummy: (c5, 0.094615ns)
signal Z2o2_normal :  std_logic_vector(10 downto 0);
   -- timing of Z2o2_normal: (c5, 0.094615ns)
signal addFinalLog1pY :  std_logic_vector(20 downto 0);
   -- timing of addFinalLog1pY: (c5, 0.644615ns)
signal Log1p_normal :  std_logic_vector(20 downto 0);
   -- timing of Log1p_normal: (c6, 0.044615ns)
signal L0 :  std_logic_vector(29 downto 0);
   -- timing of L0: (c0, 0.550000ns)
signal L0_copy28 :  std_logic_vector(29 downto 0);
   -- timing of L0_copy28: (c0, 0.000000ns)
signal S1 :  std_logic_vector(29 downto 0);
   -- timing of S1: (c0, 0.550000ns)
signal L1 :  std_logic_vector(24 downto 0);
   -- timing of L1: (c1, 1.110000ns)
signal L1_copy31 :  std_logic_vector(24 downto 0);
   -- timing of L1_copy31: (c1, 0.560000ns)
signal sopX1 :  std_logic_vector(29 downto 0);
   -- timing of sopX1: (c1, 1.110000ns)
signal S2 :  std_logic_vector(29 downto 0);
   -- timing of S2: (c2, 0.610000ns)
signal almostLog :  std_logic_vector(29 downto 0);
   -- timing of almostLog: (c2, 0.610000ns)
signal adderLogF_normalY :  std_logic_vector(29 downto 0);
   -- timing of adderLogF_normalY: (c6, 0.044615ns)
signal LogF_normal :  std_logic_vector(29 downto 0);
   -- timing of LogF_normal: (c6, 1.334615ns)
signal absELog2 :  std_logic_vector(28 downto 0);
   -- timing of absELog2: (c1, 1.650000ns)
signal absELog2_pad :  std_logic_vector(37 downto 0);
   -- timing of absELog2_pad: (c1, 1.650000ns)
signal LogF_normal_pad :  std_logic_vector(37 downto 0);
   -- timing of LogF_normal_pad: (c6, 1.334615ns)
signal lnaddX :  std_logic_vector(37 downto 0);
   -- timing of lnaddX: (c1, 1.650000ns)
signal lnaddY :  std_logic_vector(37 downto 0);
   -- timing of lnaddY: (c6, 1.334615ns)
signal Log_normal :  std_logic_vector(37 downto 0);
   -- timing of Log_normal: (c8, 0.114615ns)
signal Log_normal_normd :  std_logic_vector(29 downto 0);
   -- timing of Log_normal_normd: (c11, 0.304615ns)
signal E_normal :  std_logic_vector(4 downto 0);
   -- timing of E_normal: (c10, 1.554615ns)
signal Z2o2_small_bs :  std_logic_vector(13 downto 0);
   -- timing of Z2o2_small_bs: (c5, 0.094615ns)
signal Z2o2_small_s :  std_logic_vector(26 downto 0);
   -- timing of Z2o2_small_s: (c6, 0.102308ns)
signal Z2o2_small :  std_logic_vector(22 downto 0);
   -- timing of Z2o2_small: (c6, 0.102308ns)
signal Z_small :  std_logic_vector(22 downto 0);
   -- timing of Z_small: (c4, 1.344615ns)
signal Log_smallY :  std_logic_vector(22 downto 0);
   -- timing of Log_smallY: (c6, 0.102308ns)
signal nsRCin :  std_logic;
   -- timing of nsRCin: (c0, 0.550000ns)
signal Log_small :  std_logic_vector(22 downto 0);
   -- timing of Log_small: (c6, 1.322308ns)
signal E0_sub :  std_logic_vector(1 downto 0);
   -- timing of E0_sub: (c6, 1.322308ns)
signal ufl, ufl_d1, ufl_d2, ufl_d3, ufl_d4, ufl_d5, ufl_d6, ufl_d7, ufl_d8, ufl_d9, ufl_d10, ufl_d11 :  std_logic;
   -- timing of ufl: (c0, 0.000000ns)
signal E_small, E_small_d1, E_small_d2, E_small_d3, E_small_d4 :  std_logic_vector(7 downto 0);
   -- timing of E_small: (c6, 1.322308ns)
signal Log_small_normd, Log_small_normd_d1, Log_small_normd_d2, Log_small_normd_d3, Log_small_normd_d4, Log_small_normd_d5 :  std_logic_vector(20 downto 0);
   -- timing of Log_small_normd: (c6, 1.322308ns)
signal E0offset, E0offset_d1, E0offset_d2, E0offset_d3, E0offset_d4, E0offset_d5, E0offset_d6, E0offset_d7, E0offset_d8, E0offset_d9, E0offset_d10 :  std_logic_vector(7 downto 0);
   -- timing of E0offset: (c0, 0.000000ns)
signal ER, ER_d1 :  std_logic_vector(7 downto 0);
   -- timing of ER: (c10, 1.554615ns)
signal Log_g :  std_logic_vector(20 downto 0);
   -- timing of Log_g: (c11, 0.304615ns)
signal round :  std_logic;
   -- timing of round: (c11, 0.304615ns)
signal fraX :  std_logic_vector(24 downto 0);
   -- timing of fraX: (c11, 0.304615ns)
signal fraY :  std_logic_vector(24 downto 0);
   -- timing of fraY: (c11, 0.304615ns)
signal EFR :  std_logic_vector(24 downto 0);
   -- timing of EFR: (c11, 1.544615ns)
signal Rexn :  std_logic_vector(2 downto 0);
   -- timing of Rexn: (c11, 0.854615ns)
constant g: positive := 4;
constant log2wF: positive := 5;
constant pfinal: positive := 9;
constant sfinal: positive := 21;
constant targetprec: positive := 30;
constant wE: positive := 8;
constant wF: positive := 17;
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            XExnSgn_d1 <=  XExnSgn;
            XExnSgn_d2 <=  XExnSgn_d1;
            XExnSgn_d3 <=  XExnSgn_d2;
            XExnSgn_d4 <=  XExnSgn_d3;
            XExnSgn_d5 <=  XExnSgn_d4;
            XExnSgn_d6 <=  XExnSgn_d5;
            XExnSgn_d7 <=  XExnSgn_d6;
            XExnSgn_d8 <=  XExnSgn_d7;
            XExnSgn_d9 <=  XExnSgn_d8;
            XExnSgn_d10 <=  XExnSgn_d9;
            XExnSgn_d11 <=  XExnSgn_d10;
            Y0_d1 <=  Y0;
            sR_d1 <=  sR;
            sR_d2 <=  sR_d1;
            sR_d3 <=  sR_d2;
            sR_d4 <=  sR_d3;
            sR_d5 <=  sR_d4;
            sR_d6 <=  sR_d5;
            sR_d7 <=  sR_d6;
            sR_d8 <=  sR_d7;
            sR_d9 <=  sR_d8;
            sR_d10 <=  sR_d9;
            sR_d11 <=  sR_d10;
            EeqZero_d1 <=  EeqZero;
            EeqZero_d2 <=  EeqZero_d1;
            EeqZero_d3 <=  EeqZero_d2;
            EeqZero_d4 <=  EeqZero_d3;
            lzo_d1 <=  lzo;
            lzo_d2 <=  lzo_d1;
            lzo_d3 <=  lzo_d2;
            pfinal_s_d1 <=  pfinal_s;
            pfinal_s_d2 <=  pfinal_s_d1;
            pfinal_s_d3 <=  pfinal_s_d2;
            doRR_d1 <=  doRR;
            doRR_d2 <=  doRR_d1;
            small_d1 <=  small;
            small_d2 <=  small_d1;
            small_d3 <=  small_d2;
            small_d4 <=  small_d3;
            small_d5 <=  small_d4;
            small_d6 <=  small_d5;
            small_d7 <=  small_d6;
            small_absZ0_normd_d1 <=  small_absZ0_normd;
            InvA0_d1 <=  InvA0;
            A1_d1 <=  A1;
            ZM1_d1 <=  ZM1;
            Zfinal_d1 <=  Zfinal;
            Zfinal_d2 <=  Zfinal_d1;
            ufl_d1 <=  ufl;
            ufl_d2 <=  ufl_d1;
            ufl_d3 <=  ufl_d2;
            ufl_d4 <=  ufl_d3;
            ufl_d5 <=  ufl_d4;
            ufl_d6 <=  ufl_d5;
            ufl_d7 <=  ufl_d6;
            ufl_d8 <=  ufl_d7;
            ufl_d9 <=  ufl_d8;
            ufl_d10 <=  ufl_d9;
            ufl_d11 <=  ufl_d10;
            E_small_d1 <=  E_small;
            E_small_d2 <=  E_small_d1;
            E_small_d3 <=  E_small_d2;
            E_small_d4 <=  E_small_d3;
            Log_small_normd_d1 <=  Log_small_normd;
            Log_small_normd_d2 <=  Log_small_normd_d1;
            Log_small_normd_d3 <=  Log_small_normd_d2;
            Log_small_normd_d4 <=  Log_small_normd_d3;
            Log_small_normd_d5 <=  Log_small_normd_d4;
            E0offset_d1 <=  E0offset;
            E0offset_d2 <=  E0offset_d1;
            E0offset_d3 <=  E0offset_d2;
            E0offset_d4 <=  E0offset_d3;
            E0offset_d5 <=  E0offset_d4;
            E0offset_d6 <=  E0offset_d5;
            E0offset_d7 <=  E0offset_d6;
            E0offset_d8 <=  E0offset_d7;
            E0offset_d9 <=  E0offset_d8;
            E0offset_d10 <=  E0offset_d9;
            ER_d1 <=  ER;
         end if;
      end process;
   XExnSgn <=  X(wE+wF+2 downto wE+wF);
   FirstBit <=  X(wF-1);
   Y0 <= "1" & X(wF-1 downto 0) & "0" when FirstBit = '0' else "01" & X(wF-1 downto 0);
   Y0h <= Y0(wF downto 1);
   -- Sign of the result;
   sR <= '0'   when  (X(wE+wF-1 downto wF) = ('0' & (wE-2 downto 0 => '1')))  -- binade [1..2)
     else not X(wE+wF-1);                -- MSB of exponent
   absZ0 <=   Y0(wF-pfinal+1 downto 0)          when (sR='0') else
             ((wF-pfinal+1 downto 0 => '0') - Y0(wF-pfinal+1 downto 0));
   E <= (X(wE+wF-1 downto wF)) - ("0" & (wE-2 downto 1 => '1') & (not FirstBit));
   absE <= ((wE-1 downto 0 => '0') - E)   when sR = '1' else E;
   EeqZero <= '1' when E=(wE-1 downto 0 => '0') else '0';
   lzoc1: LZOC_17_Freq500_uid11
      port map ( clk  => clk,
                 I => Y0h,
                 OZB => FirstBit,
                 O => lzo);
   pfinal_s <= "01001";
   shiftval <= ('0' & lzo) - ('0' & pfinal_s_d3); 
   shiftvalinL <= shiftval(3 downto 0);
   shiftvalinR <= shiftval(3 downto 0);
   doRR <= shiftval(log2wF); -- sign of the result
   small <= EeqZero_d4 and not(doRR_d1);
   -- The left shifter for the 'small' case
   small_lshift: LeftShifter10_by_max_10_Freq500_uid13
      port map ( clk  => clk,
                 S => shiftvalinL,
                 X => absZ0,
                 R => small_absZ0_normd_full);
   small_absZ0_normd <= small_absZ0_normd_full(9 downto 0); -- get rid of leading zeroes
   ---------------- The range reduction box ---------------
   A0 <= X(16 downto 10);
   -- First inv table
   InvA0Table: InvA0Table_Freq500_uid15
      port map ( X => A0,
                 Y => InvA0_copy16);
   InvA0 <= InvA0_copy16; -- output copy to hold a pipeline register if needed
   P0 <= InvA0_d1 * Y0_d1;

   Z1 <= P0(19 downto 0);

   A1 <= Z1(19 downto 15);
   B1 <= Z1(14 downto 0);
   ZM1 <= Z1;
   P1 <= A1_d1*ZM1_d1;
   Y1 <= "1" & (4 downto 0 => '0') & Z1;
   EiY1 <= Y1(25 downto 5)  when A1(4) = '1'
     else  "0" & Y1(25 downto 6);
   addXIter1 <= "0" & B1 & (4 downto 0 => '0');
   addIter1_1: IntAdder_21_Freq500_uid19
      port map ( clk  => clk,
                 Cin => '0',
                 X => addXIter1,
                 Y => EiY1,
                 R => EiYPB1);
   Pp1 <= (0 downto 0 => '1') & not(P1(24 downto 5));
   addIter2_1: IntAdder_21_Freq500_uid22
      port map ( clk  => clk,
                 Cin => '1',
                 X => EiYPB1,
                 Y => Pp1,
                 R => Z2);
   Zfinal <= Z2;
   squarerIn <= Zfinal_d2(sfinal-1 downto sfinal-14) when doRR_d2='1'
                    else (small_absZ0_normd_d1 & (3 downto 0 => '0'));  
   Z2o2_full <= squarerIn*squarerIn;
   Z2o2_full_dummy <= Z2o2_full;
   Z2o2_normal <= Z2o2_full_dummy (27  downto 17);
   addFinalLog1pY <= (pfinal downto 0  => '1') & not(Z2o2_normal);
   addFinalLog1p_normalAdder: IntAdder_21_Freq500_uid25
      port map ( clk  => clk,
                 Cin => '1',
                 X => Zfinal,
                 Y => addFinalLog1pY,
                 R => Log1p_normal);

   -- Now the log tables, as late as possible
   LogTable0: LogTable0_Freq500_uid27
      port map ( X => A0,
                 Y => L0_copy28);
   L0 <= L0_copy28; -- output copy to hold a pipeline register if needed
   S1 <= L0;
   LogTable1: LogTable1_Freq500_uid30
      port map ( X => A1,
                 Y => L1_copy31);
   L1 <= L1_copy31; -- output copy to hold a pipeline register if needed
   sopX1 <= ((29 downto 25 => '0') & L1);
   adderS1: IntAdder_30_Freq500_uid34
      port map ( clk  => clk,
                 Cin => '0',
                 X => S1,
                 Y => sopX1,
                 R => S2);
   almostLog <= S2;
   adderLogF_normalY <= ((targetprec-1 downto sfinal => '0') & Log1p_normal);
   adderLogF_normal: IntAdder_30_Freq500_uid37
      port map ( clk  => clk,
                 Cin => '0',
                 X => almostLog,
                 Y => adderLogF_normalY,
                 R => LogF_normal);
   MulLog2: FixRealKCM_Freq500_uid39
      port map ( clk  => clk,
                 X => absE,
                 R => absELog2);
   absELog2_pad <=   absELog2 & (targetprec-wF-g-1 downto 0 => '0');       
   LogF_normal_pad <= (wE-1  downto 0 => LogF_normal(targetprec-1))  & LogF_normal;
   lnaddX <= absELog2_pad;
   lnaddY <= LogF_normal_pad when sR_d6='0' else not(LogF_normal_pad); 
   lnadder: IntAdder_38_Freq500_uid51
      port map ( clk  => clk,
                 Cin => sR,
                 X => lnaddX,
                 Y => lnaddY,
                 R => Log_normal);
   final_norm: Normalizer_Z_38_30_16_Freq500_uid53
      port map ( clk  => clk,
                 X => Log_normal,
                 Count => E_normal,
                 R => Log_normal_normd);
   Z2o2_small_bs <= Z2o2_full_dummy(27 downto 14);
   ao_rshift: RightShifter14_by_max_13_Freq500_uid55
      port map ( clk  => clk,
                 S => shiftvalinR,
                 X => Z2o2_small_bs,
                 R => Z2o2_small_s);
     -- send the MSB to position pfinal
   Z2o2_small <=  (pfinal-1 downto 0  => '0') & Z2o2_small_s(26 downto 13);
   -- mantissa will be either Y0-z^2/2  or  -Y0+z^2/2,  depending on sR  
   Z_small <= small_absZ0_normd & (12 downto 0 => '0');
   Log_smallY <= Z2o2_small when sR_d6='1' else not(Z2o2_small);
   nsRCin <= not ( sR );
   log_small_adder: IntAdder_23_Freq500_uid57
      port map ( clk  => clk,
                 Cin => nsRCin,
                 X => Z_small,
                 Y => Log_smallY,
                 R => Log_small);
   -- Possibly subtract 1 or 2 to the exponent, depending on the LZC of Log_small
   E0_sub <=   "11" when Log_small(wF+g+1) = '1'
          else "10" when Log_small(wF+g+1 downto wF+g) = "01"
          else "01" ;
   -- The smallest log will be log(1+2^{-wF}) \approx 2^{-wF}  = 2^-17
   -- The smallest representable number is 2^{1-2^(wE-1)} = 2^-127
   -- No underflow possible
   ufl <= '0';
   E_small <=  ("0" & (wE-2 downto 2 => '1') & E0_sub)  -  ((wE-1 downto 5 => '0') & lzo_d3) ;
   Log_small_normd <= Log_small(wF+g+1 downto 2) when Log_small(wF+g+1)='1'
           else Log_small(wF+g downto 1)  when Log_small(wF+g)='1'  -- remove the first zero
           else Log_small(wF+g-1 downto 0)  ; -- remove two zeroes (extremely rare, 001000000 only)
   E0offset <= "10000110"; -- E0 + wE 
   ER <= E_small_d4(7 downto 0) when small_d6='1'
      else E0offset_d10 - ((7 downto 5 => '0') & E_normal);
   Log_g <=  Log_small_normd_d5(wF+g-2 downto 0) & "0" when small_d7='1'           -- remove implicit 1
      else Log_normal_normd(targetprec-2 downto targetprec-wF-g-1 );  -- remove implicit 1
   round <= Log_g(g-1) ; -- sticky is always 1 for a transcendental function 
   -- if round leads to a change of binade, the carry propagation magically updates both mantissa and exponent
   fraX <= (ER_d1 & Log_g(wF+g-1 downto g)) ; 
   fraY <= ((wE+wF-1 downto 1 => '0') & round); 
   finalRoundAdder: IntAdder_25_Freq500_uid60
      port map ( clk  => clk,
                 Cin => '0',
                 X => fraX,
                 Y => fraY,
                 R => EFR);
   Rexn <= "110" when ((XExnSgn_d11(2) and (XExnSgn_d11(1) or XExnSgn_d11(0))) or (XExnSgn_d11(1) and XExnSgn_d11(0))) = '1' else
                              "101" when XExnSgn_d11(2 downto 1) = "00"  else
                              "100" when XExnSgn_d11(2 downto 1) = "10"  else
                              "00" & sR_d11 when (((Log_normal_normd(targetprec-1)='0') and (small_d7='0')) or ( (Log_small_normd_d5 (wF+g-1)='0') and (small_d7='1'))) or (ufl_d11 = '1' and small_d7='1') else
                               "01" & sR_d11;
   R<=  Rexn & EFR;
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplier_18x8_21_Freq500_uid65
-- VHDL generated for DummyFPGA @ 500MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Martin Kumm, Florent de Dinechin, Andreas Böttcher, Kinga Illyes, Bogdan Popa, Bogdan Pasca, 2012-
--------------------------------------------------------------------------------
-- Pipeline depth: 11 cycles
-- Clock period (ns): 2
-- Target frequency (MHz): 500
-- Input signals: X Y
-- Output signals: R
--  approx. input signal timings: X: (c11, 1.544615ns)Y: (c0, 0.000000ns)
--  approx. output signal timings: R: (c11, 1.544615ns)

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity IntMultiplier_18x8_21_Freq500_uid65 is
    port (clk : in std_logic;
          X : in  std_logic_vector(17 downto 0);
          Y : in  std_logic_vector(7 downto 0);
          R : out  std_logic_vector(20 downto 0)   );
end entity;

architecture arch of IntMultiplier_18x8_21_Freq500_uid65 is
signal XX_m66 :  std_logic_vector(17 downto 0);
   -- timing of XX_m66: (c11, 1.544615ns)
signal YY_m66 :  std_logic_vector(7 downto 0);
   -- timing of YY_m66: (c0, 0.000000ns)
signal XX :  unsigned(-1+18 downto 0);
   -- timing of XX: (c11, 1.544615ns)
signal YY, YY_d1, YY_d2, YY_d3, YY_d4, YY_d5, YY_d6, YY_d7, YY_d8, YY_d9, YY_d10, YY_d11 :  unsigned(-1+8 downto 0);
   -- timing of YY: (c0, 0.000000ns)
signal RR :  unsigned(-1+26 downto 0);
   -- timing of RR: (c11, 1.544615ns)
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            YY_d1 <=  YY;
            YY_d2 <=  YY_d1;
            YY_d3 <=  YY_d2;
            YY_d4 <=  YY_d3;
            YY_d5 <=  YY_d4;
            YY_d6 <=  YY_d5;
            YY_d7 <=  YY_d6;
            YY_d8 <=  YY_d7;
            YY_d9 <=  YY_d8;
            YY_d10 <=  YY_d9;
            YY_d11 <=  YY_d10;
         end if;
      end process;
   XX_m66 <= X ;
   YY_m66 <= Y ;
   XX <= unsigned(X);
   YY <= unsigned(Y);
   RR <= XX*YY_d11;
   R <= std_logic_vector(RR(25 downto 5));
end architecture;

--------------------------------------------------------------------------------
--                         IntAdder_28_Freq500_uid69
-- VHDL generated for DummyFPGA @ 500MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin (2008-2016)
--------------------------------------------------------------------------------
-- Pipeline depth: 13 cycles
-- Clock period (ns): 2
-- Target frequency (MHz): 500
-- Input signals: X Y Cin
-- Output signals: R
--  approx. input signal timings: X: (c13, 0.124615ns)Y: (c0, 0.000000ns)Cin: (c0, 0.000000ns)
--  approx. output signal timings: R: (c13, 1.394615ns)

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntAdder_28_Freq500_uid69 is
    port (clk : in std_logic;
          X : in  std_logic_vector(27 downto 0);
          Y : in  std_logic_vector(27 downto 0);
          Cin : in  std_logic;
          R : out  std_logic_vector(27 downto 0)   );
end entity;

architecture arch of IntAdder_28_Freq500_uid69 is
signal Rtmp :  std_logic_vector(27 downto 0);
   -- timing of Rtmp: (c13, 1.394615ns)
signal Y_d1, Y_d2, Y_d3, Y_d4, Y_d5, Y_d6, Y_d7, Y_d8, Y_d9, Y_d10, Y_d11, Y_d12, Y_d13 :  std_logic_vector(27 downto 0);
   -- timing of Y: (c0, 0.000000ns)
signal Cin_d1, Cin_d2, Cin_d3, Cin_d4, Cin_d5, Cin_d6, Cin_d7, Cin_d8, Cin_d9, Cin_d10, Cin_d11, Cin_d12, Cin_d13 :  std_logic;
   -- timing of Cin: (c0, 0.000000ns)
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            Y_d1 <=  Y;
            Y_d2 <=  Y_d1;
            Y_d3 <=  Y_d2;
            Y_d4 <=  Y_d3;
            Y_d5 <=  Y_d4;
            Y_d6 <=  Y_d5;
            Y_d7 <=  Y_d6;
            Y_d8 <=  Y_d7;
            Y_d9 <=  Y_d8;
            Y_d10 <=  Y_d9;
            Y_d11 <=  Y_d10;
            Y_d12 <=  Y_d11;
            Y_d13 <=  Y_d12;
            Cin_d1 <=  Cin;
            Cin_d2 <=  Cin_d1;
            Cin_d3 <=  Cin_d2;
            Cin_d4 <=  Cin_d3;
            Cin_d5 <=  Cin_d4;
            Cin_d6 <=  Cin_d5;
            Cin_d7 <=  Cin_d6;
            Cin_d8 <=  Cin_d7;
            Cin_d9 <=  Cin_d8;
            Cin_d10 <=  Cin_d9;
            Cin_d11 <=  Cin_d10;
            Cin_d12 <=  Cin_d11;
            Cin_d13 <=  Cin_d12;
         end if;
      end process;
   Rtmp <= X + Y_d13 + Cin_d13;
   R <= Rtmp;
end architecture;

--------------------------------------------------------------------------------
--                      FPMult_8_17_uid62_Freq500_uid63
-- VHDL generated for DummyFPGA @ 500MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin 2008-2021
--------------------------------------------------------------------------------
-- Pipeline depth: 13 cycles
-- Clock period (ns): 2
-- Target frequency (MHz): 500
-- Input signals: X Y
-- Output signals: R
--  approx. input signal timings: X: (c11, 1.544615ns)Y: (c0, 0.000000ns)
--  approx. output signal timings: R: (c13, 1.394615ns)

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity FPMult_8_17_uid62_Freq500_uid63 is
    port (clk : in std_logic;
          X : in  std_logic_vector(8+17+2 downto 0);
          Y : in  std_logic_vector(8+7+2 downto 0);
          R : out  std_logic_vector(8+18+2 downto 0)   );
end entity;

architecture arch of FPMult_8_17_uid62_Freq500_uid63 is
   component IntMultiplier_18x8_21_Freq500_uid65 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(17 downto 0);
             Y : in  std_logic_vector(7 downto 0);
             R : out  std_logic_vector(20 downto 0)   );
   end component;

   component IntAdder_28_Freq500_uid69 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(27 downto 0);
             Y : in  std_logic_vector(27 downto 0);
             Cin : in  std_logic;
             R : out  std_logic_vector(27 downto 0)   );
   end component;

signal sign, sign_d1, sign_d2 :  std_logic;
   -- timing of sign: (c11, 1.594615ns)
signal expX, expX_d1 :  std_logic_vector(7 downto 0);
   -- timing of expX: (c11, 1.544615ns)
signal expY, expY_d1, expY_d2, expY_d3, expY_d4, expY_d5, expY_d6, expY_d7, expY_d8, expY_d9, expY_d10, expY_d11, expY_d12 :  std_logic_vector(7 downto 0);
   -- timing of expY: (c0, 0.000000ns)
signal expSumPreSub, expSumPreSub_d1 :  std_logic_vector(9 downto 0);
   -- timing of expSumPreSub: (c12, 0.834615ns)
signal bias, bias_d1, bias_d2, bias_d3, bias_d4, bias_d5, bias_d6, bias_d7, bias_d8, bias_d9, bias_d10, bias_d11, bias_d12, bias_d13 :  std_logic_vector(9 downto 0);
   -- timing of bias: (c0, 0.000000ns)
signal expSum :  std_logic_vector(9 downto 0);
   -- timing of expSum: (c13, 0.124615ns)
signal sigX :  std_logic_vector(17 downto 0);
   -- timing of sigX: (c11, 1.544615ns)
signal sigY :  std_logic_vector(7 downto 0);
   -- timing of sigY: (c0, 0.000000ns)
signal sigProd, sigProd_d1 :  std_logic_vector(20 downto 0);
   -- timing of sigProd: (c11, 1.544615ns)
signal excSel :  std_logic_vector(3 downto 0);
   -- timing of excSel: (c11, 1.544615ns)
signal exc, exc_d1, exc_d2 :  std_logic_vector(1 downto 0);
   -- timing of exc: (c11, 1.594615ns)
signal norm, norm_d1, norm_d2 :  std_logic;
   -- timing of norm: (c11, 1.544615ns)
signal expPostNorm :  std_logic_vector(9 downto 0);
   -- timing of expPostNorm: (c13, 0.124615ns)
signal sigProdExt, sigProdExt_d1 :  std_logic_vector(20 downto 0);
   -- timing of sigProdExt: (c12, 0.294615ns)
signal expSig :  std_logic_vector(27 downto 0);
   -- timing of expSig: (c13, 0.124615ns)
signal round :  std_logic;
   -- timing of round: (c0, 0.000000ns)
signal expSigPostRound :  std_logic_vector(27 downto 0);
   -- timing of expSigPostRound: (c13, 1.394615ns)
signal excPostNorm :  std_logic_vector(1 downto 0);
   -- timing of excPostNorm: (c13, 1.394615ns)
signal finalExc :  std_logic_vector(1 downto 0);
   -- timing of finalExc: (c13, 1.394615ns)
signal Y_d1, Y_d2, Y_d3, Y_d4, Y_d5, Y_d6, Y_d7, Y_d8, Y_d9, Y_d10, Y_d11 :  std_logic_vector(8+7+2 downto 0);
   -- timing of Y: (c0, 0.000000ns)
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            sign_d1 <=  sign;
            sign_d2 <=  sign_d1;
            expX_d1 <=  expX;
            expY_d1 <=  expY;
            expY_d2 <=  expY_d1;
            expY_d3 <=  expY_d2;
            expY_d4 <=  expY_d3;
            expY_d5 <=  expY_d4;
            expY_d6 <=  expY_d5;
            expY_d7 <=  expY_d6;
            expY_d8 <=  expY_d7;
            expY_d9 <=  expY_d8;
            expY_d10 <=  expY_d9;
            expY_d11 <=  expY_d10;
            expY_d12 <=  expY_d11;
            expSumPreSub_d1 <=  expSumPreSub;
            bias_d1 <=  bias;
            bias_d2 <=  bias_d1;
            bias_d3 <=  bias_d2;
            bias_d4 <=  bias_d3;
            bias_d5 <=  bias_d4;
            bias_d6 <=  bias_d5;
            bias_d7 <=  bias_d6;
            bias_d8 <=  bias_d7;
            bias_d9 <=  bias_d8;
            bias_d10 <=  bias_d9;
            bias_d11 <=  bias_d10;
            bias_d12 <=  bias_d11;
            bias_d13 <=  bias_d12;
            sigProd_d1 <=  sigProd;
            exc_d1 <=  exc;
            exc_d2 <=  exc_d1;
            norm_d1 <=  norm;
            norm_d2 <=  norm_d1;
            sigProdExt_d1 <=  sigProdExt;
            Y_d1 <=  Y;
            Y_d2 <=  Y_d1;
            Y_d3 <=  Y_d2;
            Y_d4 <=  Y_d3;
            Y_d5 <=  Y_d4;
            Y_d6 <=  Y_d5;
            Y_d7 <=  Y_d6;
            Y_d8 <=  Y_d7;
            Y_d9 <=  Y_d8;
            Y_d10 <=  Y_d9;
            Y_d11 <=  Y_d10;
         end if;
      end process;
   sign <= X(25) xor Y_d11(15);
   expX <= X(24 downto 17);
   expY <= Y(14 downto 7);
   expSumPreSub <= ("00" & expX_d1) + ("00" & expY_d12);
   bias <= CONV_STD_LOGIC_VECTOR(127,10);
   expSum <= expSumPreSub_d1 - bias_d13;
   sigX <= "1" & X(16 downto 0);
   sigY <= "1" & Y(6 downto 0);
   SignificandMultiplication: IntMultiplier_18x8_21_Freq500_uid65
      port map ( clk  => clk,
                 X => sigX,
                 Y => sigY,
                 R => sigProd);
   excSel <= X(27 downto 26) & Y_d11(17 downto 16);
   with excSel  select  
   exc <= "00" when  "0000" | "0001" | "0100", 
          "01" when "0101",
          "10" when "0110" | "1001" | "1010" ,
          "11" when others;
   norm <= sigProd(20);
   -- exponent update
   expPostNorm <= expSum + ("000000000" & norm_d2);
   -- significand normalization shift
   sigProdExt <= sigProd_d1(19 downto 0) & "0" when norm_d1='1' else
                         sigProd_d1(18 downto 0) & "00";
   expSig <= expPostNorm & sigProdExt_d1(20 downto 3);
   round <= '1' ;
   RoundingAdder: IntAdder_28_Freq500_uid69
      port map ( clk  => clk,
                 Cin => round,
                 X => expSig,
                 Y => "0000000000000000000000000000",
                 R => expSigPostRound);
   with expSigPostRound(27 downto 26)  select 
   excPostNorm <=  "01"  when  "00",
                               "10"             when "01", 
                               "00"             when "11"|"10",
                               "11"             when others;
   with exc_d2  select  
   finalExc <= exc_d2 when  "11"|"10"|"00",
                       excPostNorm when others; 
   R <= finalExc & sign_d2 & expSigPostRound(25 downto 0);
end architecture;

--------------------------------------------------------------------------------
--                   LeftShifter19_by_max_16_Freq500_uid73
-- VHDL generated for DummyFPGA @ 500MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca (2008-2011), Florent de Dinechin (2008-2019)
--------------------------------------------------------------------------------
-- Pipeline depth: 2 cycles
-- Clock period (ns): 2
-- Target frequency (MHz): 500
-- Input signals: X S
-- Output signals: R
--  approx. input signal timings: X: (c13, 1.394615ns)S: (c14, 0.684615ns)
--  approx. output signal timings: R: (c15, 0.846154ns)

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity LeftShifter19_by_max_16_Freq500_uid73 is
    port (clk : in std_logic;
          X : in  std_logic_vector(18 downto 0);
          S : in  std_logic_vector(4 downto 0);
          R : out  std_logic_vector(34 downto 0)   );
end entity;

architecture arch of LeftShifter19_by_max_16_Freq500_uid73 is
signal ps, ps_d1 :  std_logic_vector(4 downto 0);
   -- timing of ps: (c14, 0.684615ns)
signal level0, level0_d1 :  std_logic_vector(18 downto 0);
   -- timing of level0: (c13, 1.394615ns)
signal level1 :  std_logic_vector(19 downto 0);
   -- timing of level1: (c14, 0.684615ns)
signal level2 :  std_logic_vector(21 downto 0);
   -- timing of level2: (c14, 1.573077ns)
signal level3, level3_d1 :  std_logic_vector(25 downto 0);
   -- timing of level3: (c14, 1.573077ns)
signal level4 :  std_logic_vector(33 downto 0);
   -- timing of level4: (c15, 0.846154ns)
signal level5 :  std_logic_vector(49 downto 0);
   -- timing of level5: (c15, 0.846154ns)
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            ps_d1 <=  ps;
            level0_d1 <=  level0;
            level3_d1 <=  level3;
         end if;
      end process;
   ps<= S;
   level0<= X;
   level1<= level0_d1 & (0 downto 0 => '0') when ps(0)= '1' else     (0 downto 0 => '0') & level0_d1;
   level2<= level1 & (1 downto 0 => '0') when ps(1)= '1' else     (1 downto 0 => '0') & level1;
   level3<= level2 & (3 downto 0 => '0') when ps(2)= '1' else     (3 downto 0 => '0') & level2;
   level4<= level3_d1 & (7 downto 0 => '0') when ps_d1(3)= '1' else     (7 downto 0 => '0') & level3_d1;
   level5<= level4 & (15 downto 0 => '0') when ps_d1(4)= '1' else     (15 downto 0 => '0') & level4;
   R <= level5(34 downto 0);
end architecture;

--------------------------------------------------------------------------------
--                         IntAdder_12_Freq500_uid87
-- VHDL generated for DummyFPGA @ 500MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin (2008-2016)
--------------------------------------------------------------------------------
-- Pipeline depth: 16 cycles
-- Clock period (ns): 2
-- Target frequency (MHz): 500
-- Input signals: X Y Cin
-- Output signals: R
--  approx. input signal timings: X: (c15, 1.396154ns)Y: (c15, 1.396154ns)Cin: (c0, 0.000000ns)
--  approx. output signal timings: R: (c16, 0.706154ns)

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntAdder_12_Freq500_uid87 is
    port (clk : in std_logic;
          X : in  std_logic_vector(11 downto 0);
          Y : in  std_logic_vector(11 downto 0);
          Cin : in  std_logic;
          R : out  std_logic_vector(11 downto 0)   );
end entity;

architecture arch of IntAdder_12_Freq500_uid87 is
signal Rtmp :  std_logic_vector(11 downto 0);
   -- timing of Rtmp: (c16, 0.706154ns)
signal X_d1 :  std_logic_vector(11 downto 0);
   -- timing of X: (c15, 1.396154ns)
signal Y_d1 :  std_logic_vector(11 downto 0);
   -- timing of Y: (c15, 1.396154ns)
signal Cin_d1, Cin_d2, Cin_d3, Cin_d4, Cin_d5, Cin_d6, Cin_d7, Cin_d8, Cin_d9, Cin_d10, Cin_d11, Cin_d12, Cin_d13, Cin_d14, Cin_d15, Cin_d16 :  std_logic;
   -- timing of Cin: (c0, 0.000000ns)
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            X_d1 <=  X;
            Y_d1 <=  Y;
            Cin_d1 <=  Cin;
            Cin_d2 <=  Cin_d1;
            Cin_d3 <=  Cin_d2;
            Cin_d4 <=  Cin_d3;
            Cin_d5 <=  Cin_d4;
            Cin_d6 <=  Cin_d5;
            Cin_d7 <=  Cin_d6;
            Cin_d8 <=  Cin_d7;
            Cin_d9 <=  Cin_d8;
            Cin_d10 <=  Cin_d9;
            Cin_d11 <=  Cin_d10;
            Cin_d12 <=  Cin_d11;
            Cin_d13 <=  Cin_d12;
            Cin_d14 <=  Cin_d13;
            Cin_d15 <=  Cin_d14;
            Cin_d16 <=  Cin_d15;
         end if;
      end process;
   Rtmp <= X_d1 + Y_d1 + Cin_d16;
   R <= Rtmp;
end architecture;

--------------------------------------------------------------------------------
--                          FixRealKCM_Freq500_uid77
-- VHDL generated for DummyFPGA @ 500MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin (2007-2016)
--------------------------------------------------------------------------------
-- Pipeline depth: 1 cycles
-- Clock period (ns): 2
-- Target frequency (MHz): 500
-- Input signals: X
-- Output signals: R
--  approx. input signal timings: X: (c15, 0.846154ns)
--  approx. output signal timings: R: (c16, 0.706154ns)

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity FixRealKCM_Freq500_uid77 is
    port (clk : in std_logic;
          X : in  std_logic_vector(9 downto 0);
          R : out  std_logic_vector(7 downto 0)   );
end entity;

architecture arch of FixRealKCM_Freq500_uid77 is
   component FixRealKCM_Freq500_uid77_T0_Freq500_uid80 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(11 downto 0)   );
   end component;

   component FixRealKCM_Freq500_uid77_T1_Freq500_uid83 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(6 downto 0)   );
   end component;

   component IntAdder_12_Freq500_uid87 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(11 downto 0);
             Y : in  std_logic_vector(11 downto 0);
             Cin : in  std_logic;
             R : out  std_logic_vector(11 downto 0)   );
   end component;

signal FixRealKCM_Freq500_uid77_A0 :  std_logic_vector(4 downto 0);
   -- timing of FixRealKCM_Freq500_uid77_A0: (c15, 0.846154ns)
signal FixRealKCM_Freq500_uid77_T0 :  std_logic_vector(11 downto 0);
   -- timing of FixRealKCM_Freq500_uid77_T0: (c15, 1.396154ns)
signal FixRealKCM_Freq500_uid77_T0_copy81 :  std_logic_vector(11 downto 0);
   -- timing of FixRealKCM_Freq500_uid77_T0_copy81: (c15, 0.846154ns)
signal bh78_w0_0 :  std_logic;
   -- timing of bh78_w0_0: (c15, 1.396154ns)
signal bh78_w1_0 :  std_logic;
   -- timing of bh78_w1_0: (c15, 1.396154ns)
signal bh78_w2_0 :  std_logic;
   -- timing of bh78_w2_0: (c15, 1.396154ns)
signal bh78_w3_0 :  std_logic;
   -- timing of bh78_w3_0: (c15, 1.396154ns)
signal bh78_w4_0 :  std_logic;
   -- timing of bh78_w4_0: (c15, 1.396154ns)
signal bh78_w5_0 :  std_logic;
   -- timing of bh78_w5_0: (c15, 1.396154ns)
signal bh78_w6_0 :  std_logic;
   -- timing of bh78_w6_0: (c15, 1.396154ns)
signal bh78_w7_0 :  std_logic;
   -- timing of bh78_w7_0: (c15, 1.396154ns)
signal bh78_w8_0 :  std_logic;
   -- timing of bh78_w8_0: (c15, 1.396154ns)
signal bh78_w9_0 :  std_logic;
   -- timing of bh78_w9_0: (c15, 1.396154ns)
signal bh78_w10_0 :  std_logic;
   -- timing of bh78_w10_0: (c15, 1.396154ns)
signal bh78_w11_0 :  std_logic;
   -- timing of bh78_w11_0: (c15, 1.396154ns)
signal FixRealKCM_Freq500_uid77_A1 :  std_logic_vector(4 downto 0);
   -- timing of FixRealKCM_Freq500_uid77_A1: (c15, 0.846154ns)
signal FixRealKCM_Freq500_uid77_T1 :  std_logic_vector(6 downto 0);
   -- timing of FixRealKCM_Freq500_uid77_T1: (c15, 1.396154ns)
signal FixRealKCM_Freq500_uid77_T1_copy84 :  std_logic_vector(6 downto 0);
   -- timing of FixRealKCM_Freq500_uid77_T1_copy84: (c15, 0.846154ns)
signal bh78_w0_1 :  std_logic;
   -- timing of bh78_w0_1: (c15, 1.396154ns)
signal bh78_w1_1 :  std_logic;
   -- timing of bh78_w1_1: (c15, 1.396154ns)
signal bh78_w2_1 :  std_logic;
   -- timing of bh78_w2_1: (c15, 1.396154ns)
signal bh78_w3_1 :  std_logic;
   -- timing of bh78_w3_1: (c15, 1.396154ns)
signal bh78_w4_1 :  std_logic;
   -- timing of bh78_w4_1: (c15, 1.396154ns)
signal bh78_w5_1 :  std_logic;
   -- timing of bh78_w5_1: (c15, 1.396154ns)
signal bh78_w6_1 :  std_logic;
   -- timing of bh78_w6_1: (c15, 1.396154ns)
signal bitheapFinalAdd_bh78_In0 :  std_logic_vector(11 downto 0);
   -- timing of bitheapFinalAdd_bh78_In0: (c15, 1.396154ns)
signal bitheapFinalAdd_bh78_In1 :  std_logic_vector(11 downto 0);
   -- timing of bitheapFinalAdd_bh78_In1: (c15, 1.396154ns)
signal bitheapFinalAdd_bh78_Cin :  std_logic;
   -- timing of bitheapFinalAdd_bh78_Cin: (c0, 0.000000ns)
signal bitheapFinalAdd_bh78_Out :  std_logic_vector(11 downto 0);
   -- timing of bitheapFinalAdd_bh78_Out: (c16, 0.706154ns)
signal bitheapResult_bh78 :  std_logic_vector(11 downto 0);
   -- timing of bitheapResult_bh78: (c16, 0.706154ns)
signal OutRes :  std_logic_vector(11 downto 0);
   -- timing of OutRes: (c16, 0.706154ns)
begin
-- This operator multiplies by 1/log(2)
   FixRealKCM_Freq500_uid77_A0 <= X(9 downto 5);-- input address  m=6  l=2
   FixRealKCM_Freq500_uid77_Table0: FixRealKCM_Freq500_uid77_T0_Freq500_uid80
      port map ( X => FixRealKCM_Freq500_uid77_A0,
                 Y => FixRealKCM_Freq500_uid77_T0_copy81);
   FixRealKCM_Freq500_uid77_T0 <= FixRealKCM_Freq500_uid77_T0_copy81; -- output copy to hold a pipeline register if needed
   bh78_w0_0 <= FixRealKCM_Freq500_uid77_T0(0);
   bh78_w1_0 <= FixRealKCM_Freq500_uid77_T0(1);
   bh78_w2_0 <= FixRealKCM_Freq500_uid77_T0(2);
   bh78_w3_0 <= FixRealKCM_Freq500_uid77_T0(3);
   bh78_w4_0 <= FixRealKCM_Freq500_uid77_T0(4);
   bh78_w5_0 <= FixRealKCM_Freq500_uid77_T0(5);
   bh78_w6_0 <= FixRealKCM_Freq500_uid77_T0(6);
   bh78_w7_0 <= FixRealKCM_Freq500_uid77_T0(7);
   bh78_w8_0 <= FixRealKCM_Freq500_uid77_T0(8);
   bh78_w9_0 <= FixRealKCM_Freq500_uid77_T0(9);
   bh78_w10_0 <= FixRealKCM_Freq500_uid77_T0(10);
   bh78_w11_0 <= FixRealKCM_Freq500_uid77_T0(11);
   FixRealKCM_Freq500_uid77_A1 <= X(4 downto 0);-- input address  m=1  l=-3
   FixRealKCM_Freq500_uid77_Table1: FixRealKCM_Freq500_uid77_T1_Freq500_uid83
      port map ( X => FixRealKCM_Freq500_uid77_A1,
                 Y => FixRealKCM_Freq500_uid77_T1_copy84);
   FixRealKCM_Freq500_uid77_T1 <= FixRealKCM_Freq500_uid77_T1_copy84; -- output copy to hold a pipeline register if needed
   bh78_w0_1 <= FixRealKCM_Freq500_uid77_T1(0);
   bh78_w1_1 <= FixRealKCM_Freq500_uid77_T1(1);
   bh78_w2_1 <= FixRealKCM_Freq500_uid77_T1(2);
   bh78_w3_1 <= FixRealKCM_Freq500_uid77_T1(3);
   bh78_w4_1 <= FixRealKCM_Freq500_uid77_T1(4);
   bh78_w5_1 <= FixRealKCM_Freq500_uid77_T1(5);
   bh78_w6_1 <= FixRealKCM_Freq500_uid77_T1(6);

   -- Adding the constant bits 
      -- All the constant bits are zero, nothing to add


   bitheapFinalAdd_bh78_In0 <= "" & bh78_w11_0 & bh78_w10_0 & bh78_w9_0 & bh78_w8_0 & bh78_w7_0 & bh78_w6_0 & bh78_w5_0 & bh78_w4_0 & bh78_w3_0 & bh78_w2_0 & bh78_w1_0 & bh78_w0_0;
   bitheapFinalAdd_bh78_In1 <= "0" & "0" & "0" & "0" & "0" & bh78_w6_1 & bh78_w5_1 & bh78_w4_1 & bh78_w3_1 & bh78_w2_1 & bh78_w1_1 & bh78_w0_1;
   bitheapFinalAdd_bh78_Cin <= '0';

   bitheapFinalAdd_bh78: IntAdder_12_Freq500_uid87
      port map ( clk  => clk,
                 Cin => bitheapFinalAdd_bh78_Cin,
                 X => bitheapFinalAdd_bh78_In0,
                 Y => bitheapFinalAdd_bh78_In1,
                 R => bitheapFinalAdd_bh78_Out);
   bitheapResult_bh78 <= bitheapFinalAdd_bh78_Out(11 downto 0);
   OutRes <= bitheapResult_bh78(11 downto 0);
   R <= OutRes(11 downto 4);
end architecture;

--------------------------------------------------------------------------------
--                         IntAdder_18_Freq500_uid99
-- VHDL generated for DummyFPGA @ 500MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin (2008-2016)
--------------------------------------------------------------------------------
-- Pipeline depth: 17 cycles
-- Clock period (ns): 2
-- Target frequency (MHz): 500
-- Input signals: X Y Cin
-- Output signals: R
--  approx. input signal timings: X: (c16, 1.256154ns)Y: (c16, 1.256154ns)Cin: (c0, 0.000000ns)
--  approx. output signal timings: R: (c17, 0.626154ns)

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntAdder_18_Freq500_uid99 is
    port (clk : in std_logic;
          X : in  std_logic_vector(17 downto 0);
          Y : in  std_logic_vector(17 downto 0);
          Cin : in  std_logic;
          R : out  std_logic_vector(17 downto 0)   );
end entity;

architecture arch of IntAdder_18_Freq500_uid99 is
signal Rtmp :  std_logic_vector(17 downto 0);
   -- timing of Rtmp: (c17, 0.626154ns)
signal X_d1 :  std_logic_vector(17 downto 0);
   -- timing of X: (c16, 1.256154ns)
signal Y_d1 :  std_logic_vector(17 downto 0);
   -- timing of Y: (c16, 1.256154ns)
signal Cin_d1, Cin_d2, Cin_d3, Cin_d4, Cin_d5, Cin_d6, Cin_d7, Cin_d8, Cin_d9, Cin_d10, Cin_d11, Cin_d12, Cin_d13, Cin_d14, Cin_d15, Cin_d16, Cin_d17 :  std_logic;
   -- timing of Cin: (c0, 0.000000ns)
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            X_d1 <=  X;
            Y_d1 <=  Y;
            Cin_d1 <=  Cin;
            Cin_d2 <=  Cin_d1;
            Cin_d3 <=  Cin_d2;
            Cin_d4 <=  Cin_d3;
            Cin_d5 <=  Cin_d4;
            Cin_d6 <=  Cin_d5;
            Cin_d7 <=  Cin_d6;
            Cin_d8 <=  Cin_d7;
            Cin_d9 <=  Cin_d8;
            Cin_d10 <=  Cin_d9;
            Cin_d11 <=  Cin_d10;
            Cin_d12 <=  Cin_d11;
            Cin_d13 <=  Cin_d12;
            Cin_d14 <=  Cin_d13;
            Cin_d15 <=  Cin_d14;
            Cin_d16 <=  Cin_d15;
            Cin_d17 <=  Cin_d16;
         end if;
      end process;
   Rtmp <= X_d1 + Y_d1 + Cin_d17;
   R <= Rtmp;
end architecture;

--------------------------------------------------------------------------------
--                          FixRealKCM_Freq500_uid89
-- VHDL generated for DummyFPGA @ 500MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin (2007-2016)
--------------------------------------------------------------------------------
-- Pipeline depth: 1 cycles
-- Clock period (ns): 2
-- Target frequency (MHz): 500
-- Input signals: X
-- Output signals: R
--  approx. input signal timings: X: (c16, 0.706154ns)
--  approx. output signal timings: R: (c17, 0.626154ns)

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity FixRealKCM_Freq500_uid89 is
    port (clk : in std_logic;
          X : in  std_logic_vector(7 downto 0);
          R : out  std_logic_vector(17 downto 0)   );
end entity;

architecture arch of FixRealKCM_Freq500_uid89 is
   component FixRealKCM_Freq500_uid89_T0_Freq500_uid92 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(17 downto 0)   );
   end component;

   component FixRealKCM_Freq500_uid89_T1_Freq500_uid95 is
      port ( X : in  std_logic_vector(2 downto 0);
             Y : out  std_logic_vector(12 downto 0)   );
   end component;

   component IntAdder_18_Freq500_uid99 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(17 downto 0);
             Y : in  std_logic_vector(17 downto 0);
             Cin : in  std_logic;
             R : out  std_logic_vector(17 downto 0)   );
   end component;

signal FixRealKCM_Freq500_uid89_A0 :  std_logic_vector(4 downto 0);
   -- timing of FixRealKCM_Freq500_uid89_A0: (c16, 0.706154ns)
signal FixRealKCM_Freq500_uid89_T0 :  std_logic_vector(17 downto 0);
   -- timing of FixRealKCM_Freq500_uid89_T0: (c16, 1.256154ns)
signal FixRealKCM_Freq500_uid89_T0_copy93 :  std_logic_vector(17 downto 0);
   -- timing of FixRealKCM_Freq500_uid89_T0_copy93: (c16, 0.706154ns)
signal bh90_w0_0 :  std_logic;
   -- timing of bh90_w0_0: (c16, 1.256154ns)
signal bh90_w1_0 :  std_logic;
   -- timing of bh90_w1_0: (c16, 1.256154ns)
signal bh90_w2_0 :  std_logic;
   -- timing of bh90_w2_0: (c16, 1.256154ns)
signal bh90_w3_0 :  std_logic;
   -- timing of bh90_w3_0: (c16, 1.256154ns)
signal bh90_w4_0 :  std_logic;
   -- timing of bh90_w4_0: (c16, 1.256154ns)
signal bh90_w5_0 :  std_logic;
   -- timing of bh90_w5_0: (c16, 1.256154ns)
signal bh90_w6_0 :  std_logic;
   -- timing of bh90_w6_0: (c16, 1.256154ns)
signal bh90_w7_0 :  std_logic;
   -- timing of bh90_w7_0: (c16, 1.256154ns)
signal bh90_w8_0 :  std_logic;
   -- timing of bh90_w8_0: (c16, 1.256154ns)
signal bh90_w9_0 :  std_logic;
   -- timing of bh90_w9_0: (c16, 1.256154ns)
signal bh90_w10_0 :  std_logic;
   -- timing of bh90_w10_0: (c16, 1.256154ns)
signal bh90_w11_0 :  std_logic;
   -- timing of bh90_w11_0: (c16, 1.256154ns)
signal bh90_w12_0 :  std_logic;
   -- timing of bh90_w12_0: (c16, 1.256154ns)
signal bh90_w13_0 :  std_logic;
   -- timing of bh90_w13_0: (c16, 1.256154ns)
signal bh90_w14_0 :  std_logic;
   -- timing of bh90_w14_0: (c16, 1.256154ns)
signal bh90_w15_0 :  std_logic;
   -- timing of bh90_w15_0: (c16, 1.256154ns)
signal bh90_w16_0 :  std_logic;
   -- timing of bh90_w16_0: (c16, 1.256154ns)
signal bh90_w17_0 :  std_logic;
   -- timing of bh90_w17_0: (c16, 1.256154ns)
signal FixRealKCM_Freq500_uid89_A1 :  std_logic_vector(2 downto 0);
   -- timing of FixRealKCM_Freq500_uid89_A1: (c16, 0.706154ns)
signal FixRealKCM_Freq500_uid89_T1 :  std_logic_vector(12 downto 0);
   -- timing of FixRealKCM_Freq500_uid89_T1: (c16, 1.256154ns)
signal FixRealKCM_Freq500_uid89_T1_copy96 :  std_logic_vector(12 downto 0);
   -- timing of FixRealKCM_Freq500_uid89_T1_copy96: (c16, 0.706154ns)
signal bh90_w0_1 :  std_logic;
   -- timing of bh90_w0_1: (c16, 1.256154ns)
signal bh90_w1_1 :  std_logic;
   -- timing of bh90_w1_1: (c16, 1.256154ns)
signal bh90_w2_1 :  std_logic;
   -- timing of bh90_w2_1: (c16, 1.256154ns)
signal bh90_w3_1 :  std_logic;
   -- timing of bh90_w3_1: (c16, 1.256154ns)
signal bh90_w4_1 :  std_logic;
   -- timing of bh90_w4_1: (c16, 1.256154ns)
signal bh90_w5_1 :  std_logic;
   -- timing of bh90_w5_1: (c16, 1.256154ns)
signal bh90_w6_1 :  std_logic;
   -- timing of bh90_w6_1: (c16, 1.256154ns)
signal bh90_w7_1 :  std_logic;
   -- timing of bh90_w7_1: (c16, 1.256154ns)
signal bh90_w8_1 :  std_logic;
   -- timing of bh90_w8_1: (c16, 1.256154ns)
signal bh90_w9_1 :  std_logic;
   -- timing of bh90_w9_1: (c16, 1.256154ns)
signal bh90_w10_1 :  std_logic;
   -- timing of bh90_w10_1: (c16, 1.256154ns)
signal bh90_w11_1 :  std_logic;
   -- timing of bh90_w11_1: (c16, 1.256154ns)
signal bh90_w12_1 :  std_logic;
   -- timing of bh90_w12_1: (c16, 1.256154ns)
signal bitheapFinalAdd_bh90_In0 :  std_logic_vector(17 downto 0);
   -- timing of bitheapFinalAdd_bh90_In0: (c16, 1.256154ns)
signal bitheapFinalAdd_bh90_In1 :  std_logic_vector(17 downto 0);
   -- timing of bitheapFinalAdd_bh90_In1: (c16, 1.256154ns)
signal bitheapFinalAdd_bh90_Cin :  std_logic;
   -- timing of bitheapFinalAdd_bh90_Cin: (c0, 0.000000ns)
signal bitheapFinalAdd_bh90_Out :  std_logic_vector(17 downto 0);
   -- timing of bitheapFinalAdd_bh90_Out: (c17, 0.626154ns)
signal bitheapResult_bh90 :  std_logic_vector(17 downto 0);
   -- timing of bitheapResult_bh90: (c17, 0.626154ns)
signal OutRes :  std_logic_vector(17 downto 0);
   -- timing of OutRes: (c17, 0.626154ns)
begin
-- This operator multiplies by log(2)
   FixRealKCM_Freq500_uid89_A0 <= X(7 downto 3);-- input address  m=7  l=3
   FixRealKCM_Freq500_uid89_Table0: FixRealKCM_Freq500_uid89_T0_Freq500_uid92
      port map ( X => FixRealKCM_Freq500_uid89_A0,
                 Y => FixRealKCM_Freq500_uid89_T0_copy93);
   FixRealKCM_Freq500_uid89_T0 <= FixRealKCM_Freq500_uid89_T0_copy93; -- output copy to hold a pipeline register if needed
   bh90_w0_0 <= FixRealKCM_Freq500_uid89_T0(0);
   bh90_w1_0 <= FixRealKCM_Freq500_uid89_T0(1);
   bh90_w2_0 <= FixRealKCM_Freq500_uid89_T0(2);
   bh90_w3_0 <= FixRealKCM_Freq500_uid89_T0(3);
   bh90_w4_0 <= FixRealKCM_Freq500_uid89_T0(4);
   bh90_w5_0 <= FixRealKCM_Freq500_uid89_T0(5);
   bh90_w6_0 <= FixRealKCM_Freq500_uid89_T0(6);
   bh90_w7_0 <= FixRealKCM_Freq500_uid89_T0(7);
   bh90_w8_0 <= FixRealKCM_Freq500_uid89_T0(8);
   bh90_w9_0 <= FixRealKCM_Freq500_uid89_T0(9);
   bh90_w10_0 <= FixRealKCM_Freq500_uid89_T0(10);
   bh90_w11_0 <= FixRealKCM_Freq500_uid89_T0(11);
   bh90_w12_0 <= FixRealKCM_Freq500_uid89_T0(12);
   bh90_w13_0 <= FixRealKCM_Freq500_uid89_T0(13);
   bh90_w14_0 <= FixRealKCM_Freq500_uid89_T0(14);
   bh90_w15_0 <= FixRealKCM_Freq500_uid89_T0(15);
   bh90_w16_0 <= FixRealKCM_Freq500_uid89_T0(16);
   bh90_w17_0 <= FixRealKCM_Freq500_uid89_T0(17);
   FixRealKCM_Freq500_uid89_A1 <= X(2 downto 0);-- input address  m=2  l=0
   FixRealKCM_Freq500_uid89_Table1: FixRealKCM_Freq500_uid89_T1_Freq500_uid95
      port map ( X => FixRealKCM_Freq500_uid89_A1,
                 Y => FixRealKCM_Freq500_uid89_T1_copy96);
   FixRealKCM_Freq500_uid89_T1 <= FixRealKCM_Freq500_uid89_T1_copy96; -- output copy to hold a pipeline register if needed
   bh90_w0_1 <= FixRealKCM_Freq500_uid89_T1(0);
   bh90_w1_1 <= FixRealKCM_Freq500_uid89_T1(1);
   bh90_w2_1 <= FixRealKCM_Freq500_uid89_T1(2);
   bh90_w3_1 <= FixRealKCM_Freq500_uid89_T1(3);
   bh90_w4_1 <= FixRealKCM_Freq500_uid89_T1(4);
   bh90_w5_1 <= FixRealKCM_Freq500_uid89_T1(5);
   bh90_w6_1 <= FixRealKCM_Freq500_uid89_T1(6);
   bh90_w7_1 <= FixRealKCM_Freq500_uid89_T1(7);
   bh90_w8_1 <= FixRealKCM_Freq500_uid89_T1(8);
   bh90_w9_1 <= FixRealKCM_Freq500_uid89_T1(9);
   bh90_w10_1 <= FixRealKCM_Freq500_uid89_T1(10);
   bh90_w11_1 <= FixRealKCM_Freq500_uid89_T1(11);
   bh90_w12_1 <= FixRealKCM_Freq500_uid89_T1(12);

   -- Adding the constant bits 
      -- All the constant bits are zero, nothing to add


   bitheapFinalAdd_bh90_In0 <= "" & bh90_w17_0 & bh90_w16_0 & bh90_w15_0 & bh90_w14_0 & bh90_w13_0 & bh90_w12_0 & bh90_w11_0 & bh90_w10_0 & bh90_w9_0 & bh90_w8_0 & bh90_w7_0 & bh90_w6_0 & bh90_w5_0 & bh90_w4_0 & bh90_w3_0 & bh90_w2_0 & bh90_w1_0 & bh90_w0_0;
   bitheapFinalAdd_bh90_In1 <= "0" & "0" & "0" & "0" & "0" & bh90_w12_1 & bh90_w11_1 & bh90_w10_1 & bh90_w9_1 & bh90_w8_1 & bh90_w7_1 & bh90_w6_1 & bh90_w5_1 & bh90_w4_1 & bh90_w3_1 & bh90_w2_1 & bh90_w1_1 & bh90_w0_1;
   bitheapFinalAdd_bh90_Cin <= '0';

   bitheapFinalAdd_bh90: IntAdder_18_Freq500_uid99
      port map ( clk  => clk,
                 Cin => bitheapFinalAdd_bh90_Cin,
                 X => bitheapFinalAdd_bh90_In0,
                 Y => bitheapFinalAdd_bh90_In1,
                 R => bitheapFinalAdd_bh90_Out);
   bitheapResult_bh90 <= bitheapFinalAdd_bh90_Out(17 downto 0);
   OutRes <= bitheapResult_bh90(17 downto 0);
   R <= OutRes(17 downto 0);
end architecture;

--------------------------------------------------------------------------------
--                         IntAdder_10_Freq500_uid102
-- VHDL generated for DummyFPGA @ 500MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin (2008-2016)
--------------------------------------------------------------------------------
-- Pipeline depth: 17 cycles
-- Clock period (ns): 2
-- Target frequency (MHz): 500
-- Input signals: X Y Cin
-- Output signals: R
--  approx. input signal timings: X: (c15, 1.396154ns)Y: (c17, 0.626154ns)Cin: (c0, 0.000000ns)
--  approx. output signal timings: R: (c17, 1.716154ns)

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntAdder_10_Freq500_uid102 is
    port (clk : in std_logic;
          X : in  std_logic_vector(9 downto 0);
          Y : in  std_logic_vector(9 downto 0);
          Cin : in  std_logic;
          R : out  std_logic_vector(9 downto 0)   );
end entity;

architecture arch of IntAdder_10_Freq500_uid102 is
signal Rtmp :  std_logic_vector(9 downto 0);
   -- timing of Rtmp: (c17, 1.716154ns)
signal X_d1, X_d2 :  std_logic_vector(9 downto 0);
   -- timing of X: (c15, 1.396154ns)
signal Cin_d1, Cin_d2, Cin_d3, Cin_d4, Cin_d5, Cin_d6, Cin_d7, Cin_d8, Cin_d9, Cin_d10, Cin_d11, Cin_d12, Cin_d13, Cin_d14, Cin_d15, Cin_d16, Cin_d17 :  std_logic;
   -- timing of Cin: (c0, 0.000000ns)
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            X_d1 <=  X;
            X_d2 <=  X_d1;
            Cin_d1 <=  Cin;
            Cin_d2 <=  Cin_d1;
            Cin_d3 <=  Cin_d2;
            Cin_d4 <=  Cin_d3;
            Cin_d5 <=  Cin_d4;
            Cin_d6 <=  Cin_d5;
            Cin_d7 <=  Cin_d6;
            Cin_d8 <=  Cin_d7;
            Cin_d9 <=  Cin_d8;
            Cin_d10 <=  Cin_d9;
            Cin_d11 <=  Cin_d10;
            Cin_d12 <=  Cin_d11;
            Cin_d13 <=  Cin_d12;
            Cin_d14 <=  Cin_d13;
            Cin_d15 <=  Cin_d14;
            Cin_d16 <=  Cin_d15;
            Cin_d17 <=  Cin_d16;
         end if;
      end process;
   Rtmp <= X_d2 + Y + Cin_d17;
   R <= Rtmp;
end architecture;

--------------------------------------------------------------------------------
--                           Exp_8_7_Freq500_uid75
-- VHDL generated for DummyFPGA @ 500MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: F. de Dinechin, Bogdan Pasca, Orégane Desrentes (2008-2025)
--------------------------------------------------------------------------------
-- Pipeline depth: 3 cycles
-- Clock period (ns): 2
-- Target frequency (MHz): 500
-- Input signals: ufixX_i XSign
-- Output signals: expY K
--  approx. input signal timings: ufixX_i: (c15, 0.846154ns)XSign: (c13, 1.394615ns)
--  approx. output signal timings: expY: (c0, 0.000000ns)K: (c16, 1.786154ns)

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity Exp_8_7_Freq500_uid75 is
    port (clk : in std_logic;
          ufixX_i : in  std_logic_vector(16 downto 0);
          XSign : in  std_logic;
          expY : out  std_logic_vector(12 downto 0);
          K : out  std_logic_vector(8 downto 0)   );
end entity;

architecture arch of Exp_8_7_Freq500_uid75 is
   component FixRealKCM_Freq500_uid77 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(9 downto 0);
             R : out  std_logic_vector(7 downto 0)   );
   end component;

   component FixRealKCM_Freq500_uid89 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(7 downto 0);
             R : out  std_logic_vector(17 downto 0)   );
   end component;

   component IntAdder_10_Freq500_uid102 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(9 downto 0);
             Y : in  std_logic_vector(9 downto 0);
             Cin : in  std_logic;
             R : out  std_logic_vector(9 downto 0)   );
   end component;

   component FixFunctionByTable_Freq500_uid104 is
      port ( X : in  std_logic_vector(9 downto 0);
             Y : out  std_logic_vector(12 downto 0)   );
   end component;

signal ufixX :  unsigned(6+10 downto 0);
   -- timing of ufixX: (c15, 0.846154ns)
signal xMulIn :  unsigned(6+3 downto 0);
   -- timing of xMulIn: (c15, 0.846154ns)
signal absK :  std_logic_vector(7 downto 0);
   -- timing of absK: (c16, 0.706154ns)
signal minusAbsK :  std_logic_vector(8 downto 0);
   -- timing of minusAbsK: (c16, 1.786154ns)
signal absKLog2 :  std_logic_vector(17 downto 0);
   -- timing of absKLog2: (c17, 0.626154ns)
signal subOp1 :  std_logic_vector(9 downto 0);
   -- timing of subOp1: (c15, 1.396154ns)
signal subOp2 :  std_logic_vector(9 downto 0);
   -- timing of subOp2: (c17, 0.626154ns)
signal Y :  std_logic_vector(9 downto 0);
   -- timing of Y: (c17, 1.716154ns)
signal XSign_d1, XSign_d2, XSign_d3, XSign_d4 :  std_logic;
   -- timing of XSign: (c13, 1.394615ns)
constant g: positive := 3;
constant wE: positive := 8;
constant wF: positive := 7;
constant wFIn: positive := 7;
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            XSign_d1 <=  XSign;
            XSign_d2 <=  XSign_d1;
            XSign_d3 <=  XSign_d2;
            XSign_d4 <=  XSign_d3;
         end if;
      end process;
ufixX <= unsigned(ufixX_i);
   xMulIn <= ufixX(16 downto 7); -- fix resize from (6, -10) to (6, -3)
   MulInvLog2: FixRealKCM_Freq500_uid77
      port map ( clk  => clk,
                 X => std_logic_vector(xMulIn),
                 R => absK);
   minusAbsK <= (8 downto 0 => '0') - ('0' & absK);
   K <= minusAbsK when  XSign_d3='1'   else ('0' & absK);
   MulLog2: FixRealKCM_Freq500_uid89
      port map ( clk  => clk,
                 X => absK,
                 R => absKLog2);
   subOp1 <= std_logic_vector(ufixX(9 downto 0)) when XSign_d2='0' else not (std_logic_vector(ufixX(9 downto 0)));
   subOp2 <= absKLog2(9 downto 0) when XSign_d4='1' else not (absKLog2(9 downto 0));
   theYAdder: IntAdder_10_Freq500_uid102
      port map ( clk  => clk,
                 Cin => '1',
                 X => subOp1,
                 Y => subOp2,
                 R => Y);
   -- Now compute the exp of this fixed-point value
   ExpYTable: FixFunctionByTable_Freq500_uid104
      port map ( X => Y,
                 Y => expY);
end architecture;

--------------------------------------------------------------------------------
--                         IntAdder_17_Freq500_uid107
-- VHDL generated for DummyFPGA @ 500MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin (2008-2016)
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 2
-- Target frequency (MHz): 500
-- Input signals: X Y Cin
-- Output signals: R
--  approx. input signal timings: X: (c0, 0.000000ns)Y: (c0, 0.000000ns)Cin: (c0, 0.000000ns)
--  approx. output signal timings: R: (c0, 0.000000ns)

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntAdder_17_Freq500_uid107 is
    port (clk : in std_logic;
          X : in  std_logic_vector(16 downto 0);
          Y : in  std_logic_vector(16 downto 0);
          Cin : in  std_logic;
          R : out  std_logic_vector(16 downto 0)   );
end entity;

architecture arch of IntAdder_17_Freq500_uid107 is
signal Rtmp :  std_logic_vector(16 downto 0);
   -- timing of Rtmp: (c0, 0.000000ns)
begin
   Rtmp <= X + Y + Cin;
   R <= Rtmp;
end architecture;

--------------------------------------------------------------------------------
--                          FPExp_8_7_Freq500_uid71
-- VHDL generated for DummyFPGA @ 500MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: F. de Dinechin, Bogdan Pasca, Orégane Desrentes (2008-2025)
--------------------------------------------------------------------------------
-- Pipeline depth: -13 cycles
-- Clock period (ns): 2
-- Target frequency (MHz): 500
-- Input signals: X
-- Output signals: R
--  approx. input signal timings: X: (c13, 1.394615ns)
--  approx. output signal timings: R: (c0, 0.000000ns)

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity FPExp_8_7_Freq500_uid71 is
    port (clk : in std_logic;
          X : in  std_logic_vector(8+18+2 downto 0);
          R : out  std_logic_vector(8+7+2 downto 0)   );
end entity;

architecture arch of FPExp_8_7_Freq500_uid71 is
   component LeftShifter19_by_max_16_Freq500_uid73 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(18 downto 0);
             S : in  std_logic_vector(4 downto 0);
             R : out  std_logic_vector(34 downto 0)   );
   end component;

   component Exp_8_7_Freq500_uid75 is
      port ( clk : in std_logic;
             ufixX_i : in  std_logic_vector(16 downto 0);
             XSign : in  std_logic;
             expY : out  std_logic_vector(12 downto 0);
             K : out  std_logic_vector(8 downto 0)   );
   end component;

   component IntAdder_17_Freq500_uid107 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(16 downto 0);
             Y : in  std_logic_vector(16 downto 0);
             Cin : in  std_logic;
             R : out  std_logic_vector(16 downto 0)   );
   end component;

signal Xexn, Xexn_d1, Xexn_d2 :  std_logic_vector(1 downto 0);
   -- timing of Xexn: (c13, 1.394615ns)
signal XSign, XSign_d1, XSign_d2 :  std_logic;
   -- timing of XSign: (c13, 1.394615ns)
signal XexpField, XexpField_d1 :  std_logic_vector(7 downto 0);
   -- timing of XexpField: (c13, 1.394615ns)
signal Xfrac :  unsigned(-1+18 downto 0);
   -- timing of Xfrac: (c13, 1.394615ns)
signal e0, e0_d1, e0_d2, e0_d3, e0_d4, e0_d5, e0_d6, e0_d7, e0_d8, e0_d9, e0_d10, e0_d11, e0_d12, e0_d13, e0_d14 :  std_logic_vector(9 downto 0);
   -- timing of e0: (c0, 0.000000ns)
signal shiftVal :  std_logic_vector(9 downto 0);
   -- timing of shiftVal: (c14, 0.684615ns)
signal resultWillBeOne, resultWillBeOne_d1 :  std_logic;
   -- timing of resultWillBeOne: (c14, 0.684615ns)
signal mXu :  unsigned(0+18 downto 0);
   -- timing of mXu: (c13, 1.394615ns)
signal maxShift, maxShift_d1, maxShift_d2, maxShift_d3, maxShift_d4, maxShift_d5, maxShift_d6, maxShift_d7, maxShift_d8, maxShift_d9, maxShift_d10, maxShift_d11, maxShift_d12, maxShift_d13, maxShift_d14 :  std_logic_vector(8 downto 0);
   -- timing of maxShift: (c0, 0.000000ns)
signal overflow0, overflow0_d1 :  std_logic;
   -- timing of overflow0: (c14, 1.764615ns)
signal shiftValIn :  std_logic_vector(4 downto 0);
   -- timing of shiftValIn: (c14, 0.684615ns)
signal fixX0 :  std_logic_vector(34 downto 0);
   -- timing of fixX0: (c15, 0.846154ns)
signal ufixX :  unsigned(6+10 downto 0);
   -- timing of ufixX: (c15, 0.846154ns)
signal expY :  std_logic_vector(12 downto 0);
   -- timing of expY: (c0, 0.000000ns)
signal K :  std_logic_vector(8 downto 0);
   -- timing of K: (c16, 1.786154ns)
signal needNoNorm :  std_logic;
   -- timing of needNoNorm: (c0, 0.000000ns)
signal preRoundBiasSig :  std_logic_vector(16 downto 0);
   -- timing of preRoundBiasSig: (c0, 0.000000ns)
signal roundBit :  std_logic;
   -- timing of roundBit: (c0, 0.000000ns)
signal roundNormAddend :  std_logic_vector(16 downto 0);
   -- timing of roundNormAddend: (c0, 0.000000ns)
signal roundedExpSigRes :  std_logic_vector(16 downto 0);
   -- timing of roundedExpSigRes: (c0, 0.000000ns)
signal roundedExpSig :  std_logic_vector(16 downto 0);
   -- timing of roundedExpSig: (c0, 0.000000ns)
signal ofl1 :  std_logic;
   -- timing of ofl1: (c15, 0.514615ns)
signal ofl2 :  std_logic;
   -- timing of ofl2: (c0, 0.000000ns)
signal ofl3 :  std_logic;
   -- timing of ofl3: (c13, 1.394615ns)
signal ofl :  std_logic;
   -- timing of ofl: (c0, 0.000000ns)
signal ufl1 :  std_logic;
   -- timing of ufl1: (c0, 0.000000ns)
signal ufl2 :  std_logic;
   -- timing of ufl2: (c13, 1.394615ns)
signal ufl3 :  std_logic;
   -- timing of ufl3: (c14, 1.764615ns)
signal ufl :  std_logic;
   -- timing of ufl: (c0, 0.000000ns)
signal Rexn :  std_logic_vector(1 downto 0);
   -- timing of Rexn: (c0, 0.000000ns)
constant g: positive := 3;
constant wE: positive := 8;
constant wF: positive := 7;
constant wFIn: positive := 18;
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            Xexn_d1 <=  Xexn;
            Xexn_d2 <=  Xexn_d1;
            XSign_d1 <=  XSign;
            XSign_d2 <=  XSign_d1;
            XexpField_d1 <=  XexpField;
            e0_d1 <=  e0;
            e0_d2 <=  e0_d1;
            e0_d3 <=  e0_d2;
            e0_d4 <=  e0_d3;
            e0_d5 <=  e0_d4;
            e0_d6 <=  e0_d5;
            e0_d7 <=  e0_d6;
            e0_d8 <=  e0_d7;
            e0_d9 <=  e0_d8;
            e0_d10 <=  e0_d9;
            e0_d11 <=  e0_d10;
            e0_d12 <=  e0_d11;
            e0_d13 <=  e0_d12;
            e0_d14 <=  e0_d13;
            resultWillBeOne_d1 <=  resultWillBeOne;
            maxShift_d1 <=  maxShift;
            maxShift_d2 <=  maxShift_d1;
            maxShift_d3 <=  maxShift_d2;
            maxShift_d4 <=  maxShift_d3;
            maxShift_d5 <=  maxShift_d4;
            maxShift_d6 <=  maxShift_d5;
            maxShift_d7 <=  maxShift_d6;
            maxShift_d8 <=  maxShift_d7;
            maxShift_d9 <=  maxShift_d8;
            maxShift_d10 <=  maxShift_d9;
            maxShift_d11 <=  maxShift_d10;
            maxShift_d12 <=  maxShift_d11;
            maxShift_d13 <=  maxShift_d12;
            maxShift_d14 <=  maxShift_d13;
            overflow0_d1 <=  overflow0;
         end if;
      end process;
   Xexn <= X(wE+wFIn+2 downto wE+wFIn+1);
   XSign <= X(wE+wFIn);
   XexpField <= X(wE+wFIn-1 downto wFIn);
   Xfrac <= unsigned(X(wFIn-1 downto 0));
   e0 <= conv_std_logic_vector(117, wE+2);  -- bias - (wF+g)
   shiftVal <= ("00" & XexpField_d1) - e0_d14; -- for a left shift
   -- underflow when input is shifted to zero (shiftval<0), in which case exp = 1
   resultWillBeOne <= shiftVal(wE+1);
   --  mantissa with implicit bit
   mXu <= "1" & Xfrac;
   -- Partial overflow detection
   maxShift <= conv_std_logic_vector(16, wE+1);  -- wE-2 + wF+g
   overflow0 <= not shiftVal(wE+1) when shiftVal(wE downto 0) > maxShift_d14 else '0';
   shiftValIn <= shiftVal(4 downto 0);
   mantissa_shift: LeftShifter19_by_max_16_Freq500_uid73
      port map ( clk  => clk,
                 S => shiftValIn,
                 X => std_logic_vector(mXu),
                 R => fixX0);
   ufixX <=  unsigned(fixX0(34 downto 18)) when resultWillBeOne_d1='0' else "00000000000000000";
   exp_helper: Exp_8_7_Freq500_uid75
      port map ( clk  => clk,
                 XSign => XSign,
                 ufixX_i => std_logic_vector(ufixX),
                 K => K,
                 expY => expY);
   needNoNorm <= expY(12);
   -- Rounding: all this should consume one row of LUTs
   preRoundBiasSig <= conv_std_logic_vector(127, wE+2)  & expY(11 downto 5) when needNoNorm = '1'
      else conv_std_logic_vector(126, wE+2)  & expY(10 downto 4) ;
   roundBit <= expY(4)  when needNoNorm = '1'    else expY(3) ;
   roundNormAddend <= K(8) & K & (6 downto 1 => '0') & roundBit;
   roundedExpSigOperandAdder: IntAdder_17_Freq500_uid107
      port map ( clk  => clk,
                 Cin => '0',
                 X => preRoundBiasSig,
                 Y => roundNormAddend,
                 R => roundedExpSigRes);
   roundedExpSig <= roundedExpSigRes when Xexn="01" else  "000" & (wE-2 downto 0 => '1') & (wF-1 downto 0 => '0');
   ofl1 <= not XSign_d2 and overflow0_d1 and (not Xexn_d2(1) and Xexn_d2(0)); -- input positive, normal,  very large
   ofl2 <= not XSign and (roundedExpSig(wE+wF) and not roundedExpSig(wE+wF+1)) and (not Xexn(1) and Xexn(0)); -- input positive, normal, overflowed
   ofl3 <= not XSign and Xexn(1) and not Xexn(0);  -- input was -infty
   ofl <= ofl1 or ofl2 or ofl3;
   ufl1 <= (roundedExpSig(wE+wF) and roundedExpSig(wE+wF+1))  and (not Xexn(1) and Xexn(0)); -- input normal
   ufl2 <= XSign and Xexn(1) and not Xexn(0);  -- input was -infty
   ufl3 <= XSign_d1 and overflow0  and (not Xexn_d1(1) and Xexn_d1(0)); -- input negative, normal,  very large
   ufl <= ufl1 or ufl2 or ufl3;
   Rexn <= "11" when Xexn = "11"
      else "10" when ofl='1'
      else "00" when ufl='1'
      else "01";
   R <= Rexn & '0' & roundedExpSig(14 downto 0);
end architecture;

--------------------------------------------------------------------------------
--                                 top_module
--                          (FPPow_8_7_Freq500_uid2)
-- VHDL generated for DummyFPGA @ 500MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: F. de Dinechin, C. Klein  (2008)
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 2
-- Target frequency (MHz): 500
-- Input signals: X Y
-- Output signals: R
--  approx. input signal timings: X: (c0, 0.000000ns)Y: (c0, 0.000000ns)
--  approx. output signal timings: R: (c0, 0.000000ns)

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity top_module is
    port (clk : in std_logic;
          X : in  std_logic_vector(8+7+2 downto 0);
          Y : in  std_logic_vector(8+7+2 downto 0);
          R : out  std_logic_vector(8+7+2 downto 0)   );
end entity;

architecture arch of top_module is
   component IntAdder_16_Freq500_uid5 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(15 downto 0);
             Y : in  std_logic_vector(15 downto 0);
             Cin : in  std_logic;
             R : out  std_logic_vector(15 downto 0)   );
   end component;

   component LZC_7_Freq500_uid7 is
      port ( clk : in std_logic;
             I : in  std_logic_vector(6 downto 0);
             O : out  std_logic_vector(2 downto 0)   );
   end component;

   component FPLogIterative_8_17_0_500_Freq500_uid9 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(8+17+2 downto 0);
             R : out  std_logic_vector(8+17+2 downto 0)   );
   end component;

   component FPMult_8_17_uid62_Freq500_uid63 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(8+17+2 downto 0);
             Y : in  std_logic_vector(8+7+2 downto 0);
             R : out  std_logic_vector(8+18+2 downto 0)   );
   end component;

   component FPExp_8_7_Freq500_uid71 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(8+18+2 downto 0);
             R : out  std_logic_vector(8+7+2 downto 0)   );
   end component;

signal flagsX :  std_logic_vector(1 downto 0);
   -- timing of flagsX: (c0, 0.000000ns)
signal signX, signX_d1 :  std_logic;
   -- timing of signX: (c0, 0.000000ns)
signal expFieldX :  std_logic_vector(7 downto 0);
   -- timing of expFieldX: (c0, 0.000000ns)
signal fracX :  std_logic_vector(6 downto 0);
   -- timing of fracX: (c0, 0.000000ns)
signal flagsY :  std_logic_vector(1 downto 0);
   -- timing of flagsY: (c0, 0.000000ns)
signal signY, signY_d1, signY_d2 :  std_logic;
   -- timing of signY: (c0, 0.000000ns)
signal expFieldY :  std_logic_vector(7 downto 0);
   -- timing of expFieldY: (c0, 0.000000ns)
signal fracY :  std_logic_vector(6 downto 0);
   -- timing of fracY: (c0, 0.000000ns)
signal zeroX, zeroX_d1, zeroX_d2 :  std_logic;
   -- timing of zeroX: (c0, 0.550000ns)
signal zeroY, zeroY_d1 :  std_logic;
   -- timing of zeroY: (c0, 0.550000ns)
signal normalX, normalX_d1 :  std_logic;
   -- timing of normalX: (c0, 0.550000ns)
signal normalY, normalY_d1, normalY_d2 :  std_logic;
   -- timing of normalY: (c0, 0.550000ns)
signal infX, infX_d1, infX_d2 :  std_logic;
   -- timing of infX: (c0, 0.550000ns)
signal infY, infY_d1, infY_d2 :  std_logic;
   -- timing of infY: (c0, 0.550000ns)
signal s_nan_in, s_nan_in_d1 :  std_logic;
   -- timing of s_nan_in: (c0, 0.550000ns)
signal OneExpFrac :  std_logic_vector(14 downto 0);
   -- timing of OneExpFrac: (c0, 0.000000ns)
signal ExpFracX :  std_logic_vector(15 downto 0);
   -- timing of ExpFracX: (c0, 0.000000ns)
signal OneExpFracCompl :  std_logic_vector(15 downto 0);
   -- timing of OneExpFracCompl: (c0, 0.000000ns)
signal cmpXOneRes :  std_logic_vector(15 downto 0);
   -- timing of cmpXOneRes: (c0, 1.150000ns)
signal XisOneAndNormal :  std_logic;
   -- timing of XisOneAndNormal: (c0, 0.550000ns)
signal absXgtOneAndNormal, absXgtOneAndNormal_d1, absXgtOneAndNormal_d2 :  std_logic;
   -- timing of absXgtOneAndNormal: (c0, 1.700000ns)
signal absXltOneAndNormal, absXltOneAndNormal_d1, absXltOneAndNormal_d2 :  std_logic;
   -- timing of absXltOneAndNormal: (c0, 1.700000ns)
signal fracYreverted :  std_logic_vector(6 downto 0);
   -- timing of fracYreverted: (c0, 0.000000ns)
signal Z_rightY, Z_rightY_d1 :  std_logic_vector(2 downto 0);
   -- timing of Z_rightY: (c0, 1.660000ns)
signal WeightLSBYpre, WeightLSBYpre_d1 :  std_logic_vector(8 downto 0);
   -- timing of WeightLSBYpre: (c0, 1.080000ns)
signal WeightLSBY, WeightLSBY_d1 :  std_logic_vector(8 downto 0);
   -- timing of WeightLSBY: (c1, 0.940000ns)
signal oddIntY, oddIntY_d1 :  std_logic;
   -- timing of oddIntY: (c1, 1.490000ns)
signal evenIntY :  std_logic;
   -- timing of evenIntY: (c2, 0.240000ns)
signal notIntNormalY :  std_logic;
   -- timing of notIntNormalY: (c1, 1.490000ns)
signal RisInfSpecialCase :  std_logic;
   -- timing of RisInfSpecialCase: (c2, 0.790000ns)
signal RisZeroSpecialCase :  std_logic;
   -- timing of RisZeroSpecialCase: (c2, 0.790000ns)
signal RisOne :  std_logic;
   -- timing of RisOne: (c0, 1.100000ns)
signal RisNaN :  std_logic;
   -- timing of RisNaN: (c1, 1.490000ns)
signal signR :  std_logic;
   -- timing of signR: (c1, 1.490000ns)
signal logIn :  std_logic_vector(27 downto 0);
   -- timing of logIn: (c0, 0.000000ns)
signal lnX :  std_logic_vector(8+17+2 downto 0);
   -- timing of lnX: (c11, 1.544615ns)
signal P :  std_logic_vector(8+18+2 downto 0);
   -- timing of P: (c13, 1.394615ns)
signal E :  std_logic_vector(8+7+2 downto 0);
   -- timing of E: (c0, 0.000000ns)
signal flagsE :  std_logic_vector(1 downto 0);
   -- timing of flagsE: (c0, 0.000000ns)
signal RisZeroFromExp :  std_logic;
   -- timing of RisZeroFromExp: (c0, 0.000000ns)
signal RisZero :  std_logic;
   -- timing of RisZero: (c0, 0.000000ns)
signal RisInfFromExp :  std_logic;
   -- timing of RisInfFromExp: (c0, 0.000000ns)
signal RisInf :  std_logic;
   -- timing of RisInf: (c0, 0.000000ns)
signal flagR :  std_logic_vector(1 downto 0);
   -- timing of flagR: (c0, 0.000000ns)
signal R_expfrac :  std_logic_vector(14 downto 0);
   -- timing of R_expfrac: (c0, 0.000000ns)
constant wE: positive := 8;
constant wF: positive := 7;
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            signX_d1 <=  signX;
            signY_d1 <=  signY;
            signY_d2 <=  signY_d1;
            zeroX_d1 <=  zeroX;
            zeroX_d2 <=  zeroX_d1;
            zeroY_d1 <=  zeroY;
            normalX_d1 <=  normalX;
            normalY_d1 <=  normalY;
            normalY_d2 <=  normalY_d1;
            infX_d1 <=  infX;
            infX_d2 <=  infX_d1;
            infY_d1 <=  infY;
            infY_d2 <=  infY_d1;
            s_nan_in_d1 <=  s_nan_in;
            absXgtOneAndNormal_d1 <=  absXgtOneAndNormal;
            absXgtOneAndNormal_d2 <=  absXgtOneAndNormal_d1;
            absXltOneAndNormal_d1 <=  absXltOneAndNormal;
            absXltOneAndNormal_d2 <=  absXltOneAndNormal_d1;
            Z_rightY_d1 <=  Z_rightY;
            WeightLSBYpre_d1 <=  WeightLSBYpre;
            WeightLSBY_d1 <=  WeightLSBY;
            oddIntY_d1 <=  oddIntY;
         end if;
      end process;
   flagsX <= X(wE+wF+2 downto wE+wF+1);
   signX <= X(wE+wF);
   expFieldX <= X(wE+wF-1 downto wF);
   fracX <= X(wF-1 downto 0);
   flagsY <= Y(wE+wF+2 downto wE+wF+1);
   signY <= Y(wE+wF);
   expFieldY <= Y(wE+wF-1 downto wF);
   fracY <= Y(wF-1 downto 0);
-- Inputs analysis  --
-- zero inputs--
   zeroX <= '1' when flagsX="00" else '0';
   zeroY <= '1' when flagsY="00" else '0';
-- normal inputs--
   normalX <= '1' when flagsX="01" else '0';
   normalY <= '1' when flagsY="01" else '0';
-- inf input --
   infX <= '1' when flagsX="10" else '0';
   infY <= '1' when flagsY="10" else '0';
-- NaN inputs  --
   s_nan_in <= '1' when flagsX="11" or flagsY="11" else '0';
-- Comparison of X to 1   --
   OneExpFrac <=  "0" & (6 downto 0 => '1') & (6 downto 0 => '0');
   ExpFracX<= "0" & expFieldX & fracX;
   OneExpFracCompl<=  "1" & (not OneExpFrac);
   cmpXOne: IntAdder_16_Freq500_uid5
      port map ( clk  => clk,
                 Cin => '1',
                 X => ExpFracX,
                 Y => OneExpFracCompl,
                 R => cmpXOneRes);
   XisOneAndNormal <= '1' when X = ("010" & OneExpFrac) else '0';
   absXgtOneAndNormal <= normalX and (not XisOneAndNormal) and (not cmpXOneRes(15));
   absXltOneAndNormal <= normalX and cmpXOneRes(15);
   fracYreverted <= fracY(0)&fracY(1)&fracY(2)&fracY(3)&fracY(4)&fracY(5)&fracY(6);
   FPPow_8_7_Freq500_uid2right1counter: LZC_7_Freq500_uid7
      port map ( clk  => clk,
                 I => fracYreverted,
                 O => Z_rightY);
-- compute the weight of the less significant one of the mantissa
   WeightLSBYpre <= ('0' & expFieldY)- CONV_STD_LOGIC_VECTOR(134,9);
   WeightLSBY <= WeightLSBYpre_d1 + Z_rightY_d1;
   oddIntY <= normalY_d1 when WeightLSBY = CONV_STD_LOGIC_VECTOR(0, 9) else '0'; -- LSB has null weight
   evenIntY <= normalY_d2 when WeightLSBY_d1(wE)='0' and oddIntY_d1='0' else '0'; --LSB has strictly positive weight 
   notIntNormalY <= normalY_d1 when WeightLSBY(wE)='1' else '0'; -- LSB has negative weight

-- Pow Exceptions  --
   RisInfSpecialCase  <= 
         (zeroX_d2  and  (oddIntY_d1 or evenIntY)  and signY_d2)  -- (+/- 0) ^ (negative int y)
      or (zeroX_d2 and infY_d2 and signY_d2)                      -- (+/- 0) ^ (-inf)
      or (absXgtOneAndNormal_d2   and  infY_d2  and not signY_d2) -- (|x|>1) ^ (+inf)
      or (absXltOneAndNormal_d2   and  infY_d2  and signY_d2)     -- (|x|<1) ^ (-inf)
      or (infX_d2 and  normalY_d2  and not signY_d2) ;            -- (inf) ^ (y>0)
   RisZeroSpecialCase <= 
         (zeroX_d2 and  (oddIntY_d1 or evenIntY)  and not signY_d2)  -- (+/- 0) ^ (positive int y)
      or (zeroX_d2 and  infY_d2  and not signY_d2)                   -- (+/- 0) ^ (+inf)
      or (absXltOneAndNormal_d2   and  infY_d2  and not signY_d2)    -- (|x|<1) ^ (+inf)
      or (absXgtOneAndNormal_d2   and  infY_d2  and signY_d2)        -- (|x|>1) ^ (-inf)
      or (infX_d2 and  normalY_d2  and signY_d2) ;                   -- (inf) ^ (y<0)
   RisOne <= 
         zeroY                                          -- x^0 = 1 without exception
      or (XisOneAndNormal and signX and infY)           -- (-1) ^ (-/-inf)
      or (XisOneAndNormal  and not signX);              -- (+1) ^ (whatever)
   RisNaN <= (s_nan_in_d1 and not zeroY_d1) or (normalX_d1 and signX_d1 and notIntNormalY);
   signR <= signX_d1 and (oddIntY);
   logIn <= flagsX & "0" & expFieldX & fracX & (9 downto 0 => '0') ;
   FPPow_8_7_Freq500_uid2log: FPLogIterative_8_17_0_500_Freq500_uid9
      port map ( clk  => clk,
                 X => logIn,
                 R => lnX);
   FPPow_8_7_Freq500_uid2mult: FPMult_8_17_uid62_Freq500_uid63
      port map ( clk  => clk,
                 X => lnX,
                 Y => Y,
                 R => P);
   FPPow_8_7_Freq500_uid2exp: FPExp_8_7_Freq500_uid71
      port map ( clk  => clk,
                 X => P,
                 R => E);
   flagsE <= E(wE+wF+2 downto wE+wF+1);
   RisZeroFromExp <= '1' when flagsE="00" else '0';
   RisZero <= RisZeroSpecialCase or RisZeroFromExp;
   RisInfFromExp  <= '1' when flagsE="10" else '0';
   RisInf  <= RisInfSpecialCase or RisInfFromExp;
   flagR <= 
           "11" when RisNaN='1'
      else "00" when RisZero='1'
      else "10" when RisInf='1'
      else "01";
   R_expfrac <= CONV_STD_LOGIC_VECTOR(127,8) &  CONV_STD_LOGIC_VECTOR(0, 7) when RisOne='1'
       else E(14 downto 0);
   R <= flagR & signR & R_expfrac;
end architecture;

--------------------------------------------------------------------------------
--                    TestBench_top_module_Freq500_uid109
-- VHDL generated for DummyFPGA @ 500MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Cristian Klein, Nicolas Brunie (2007-2010)
--------------------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity TestBench_top_module_Freq500_uid109 is
end entity;

architecture behavorial of TestBench_top_module_Freq500_uid109 is
   component top_module is
      port ( clk : in std_logic;
             X : in  std_logic_vector(8+7+2 downto 0);
             Y : in  std_logic_vector(8+7+2 downto 0);
             R : out  std_logic_vector(8+7+2 downto 0)   );
   end component;
signal X :  std_logic_vector(17 downto 0);
   -- timing of X: (c0, 0.000000ns)
signal Y :  std_logic_vector(17 downto 0);
   -- timing of Y: (c0, 0.000000ns)
signal R :  std_logic_vector(17 downto 0);
   -- timing of R: (c0, 0.000000ns)
signal clk :  std_logic;
   -- timing of clk: (c0, 0.000000ns)
signal rst :  std_logic;
   -- timing of rst: (c0, 0.000000ns)

 -- converts std_logic into a character
   function chr(sl: std_logic) return character is
      variable c: character;
   begin
      case sl is
         when 'U' => c:= 'U';
         when 'X' => c:= 'X';
         when '0' => c:= '0';
         when '1' => c:= '1';
         when 'Z' => c:= 'Z';
         when 'W' => c:= 'W';
         when 'L' => c:= 'L';
         when 'H' => c:= 'H';
         when '-' => c:= '-';
      end case;
      return c;
   end chr;

   -- converts bit to std_logic (1 to 1)
   function to_stdlogic(b : bit) return std_logic is
       variable sl : std_logic;
   begin
      case b is 
         when '0' => sl := '0';
         when '1' => sl := '1';
      end case;
      return sl;
   end to_stdlogic;

   -- converts std_logic into a string (1 to 1)
   function str(sl: std_logic) return string is
    variable s: string(1 to 1);
    begin
      s(1) := chr(sl);
      return s;
   end str;

   -- converts std_logic_vector into a string (binary base)
   -- (this also takes care of the fact that the range of
   --  a string is natural while a std_logic_vector may
   --  have an integer range)
   function str(slv: std_logic_vector) return string is
      variable result : string (1 to slv'length);
      variable r : integer;
   begin
      r := 1;
      for i in slv'range loop
         result(r) := chr(slv(i));
         r := r + 1;
      end loop;
      return result;
   end str;

   -- FP compare function (found vs. real)
   function fp_equal(a : std_logic_vector; b : std_logic_vector) return boolean is
   begin
      if b(b'high downto b'high-1) = "01" then
         return a = b;
      elsif b(b'high downto b'high-1) = "11" then
         return (a(a'high downto a'high-1)=b(b'high downto b'high-1));
      else
         return a(a'high downto a'high-2) = b(b'high downto b'high-2);
      end if;
   end;

   function fp_inf_or_equal(a : std_logic_vector; b : std_logic_vector) return boolean is
   begin
      if (b(b'high downto b'high-1) = "11") or (a(a'high downto a'high-1) = "11")  then
         return false; -- NaN always compare false
      else return true; -- TODO
      end if;
   end;

   -- FP subtypes for casting
   subtype fp18 is std_logic_vector(17 downto 0);
   function testLine(testCounter:integer; expectedOutputS: string(1 to 10000); expectedOutputSize: integer; R:  std_logic_vector(8+7+2 downto 0)) return boolean is
      variable expectedOutput: line;
      variable possibilityNumber : integer;
      variable testSuccess: boolean;
      variable errorMessage: string(1 to 10000);
      variable testSuccess_R: boolean;
      variable expected_R: bit_vector (17 downto 0); -- for list of values
      variable inf_R: bit_vector (17 downto 0); -- for intervals
      variable sup_R: bit_vector (17 downto 0); -- for intervals
   begin
      write(expectedOutput, expectedOutputS);
      read(expectedOutput, possibilityNumber); -- for R
      if possibilityNumber = 0 then
         -- TODO define what it means to have 0 possible output. Currently it means a test fails...
      end if;
      if possibilityNumber > 0 then -- a list of values
      testSuccess_R := false;
         for i in 1 to possibilityNumber loop
            read(expectedOutput, expected_R);
            if fp_equal(R, to_stdlogicvector(expected_R)) then
               testSuccess_R := true;
            end if;
            end loop;
      end if;
      if possibilityNumber < 0  then -- an interval
         read(expectedOutput, inf_R);
         read(expectedOutput, sup_R);
         if possibilityNumber =-1  then -- an unsigned interval
            testSuccess_R := (R >= to_stdlogicvector(inf_R)) and (R <= to_stdlogicvector(sup_R));
         elsif possibilityNumber =-2  then -- a signed interval
            testSuccess_R := (signed(R) >= signed(to_stdlogicvector(inf_R))) and (signed(R) <= signed(to_stdlogicvector(sup_R)));
         elsif possibilityNumber =-4  then -- a floating-point interval
            testSuccess_R := fp_inf_or_equal(to_stdlogicvector(inf_R), R) and fp_inf_or_equal(R, to_stdlogicvector(sup_R));
         end if;
      end if;
      if testSuccess_R = false then
         report("Test #" & integer'image(testCounter) & ", incorrect output for R: " & lf & " expected values: " & expectedOutputS(1 to expectedOutputSize) & lf  & "          result:    " & str(R) ) severity error;
      end if;
      
      testSuccess := true and testSuccess_R;
      return testSuccess;
   end testLine;

begin
   -- Ticking clock signal
   process
   begin
      clk <= '0';
      wait for 5 ns;
      clk <= '1';
      wait for 5 ns;
   end process;

   test: top_module
      port map ( clk  => clk,
                 X => X,
                 Y => Y,
                 R => R);
   -- Process that sets the inputs  (read from a file) 
   process
      variable input, expectedOutput : line; 
      variable tmpChar : character;
      file inputsFile : text is "test.input"; 
      variable V_X : bit_vector(17 downto 0);
      variable V_Y : bit_vector(17 downto 0);
      variable V_R : bit_vector(17 downto 0);
   begin
      -- Send reset
      rst <= '1';
      wait for 10 ns;
      rst <= '0';
      readline(inputsFile, input); -- skip the first line of advertising
      while not endfile(inputsFile) loop
         readline(inputsFile, input); -- skip the comment line
         readline(inputsFile, input);
         readline(inputsFile, expectedOutput); -- comment line, unused in this process
         readline(inputsFile, expectedOutput); -- unused in this process
         read(input ,V_X);
         read(input,tmpChar);
         X <= to_stdlogicvector(V_X);
         read(input ,V_Y);
         read(input,tmpChar);
         Y <= to_stdlogicvector(V_Y);
         wait for 10 ns;
      end loop;
         wait for 100 ns; -- wait for pipeline to flush (and some more)
   end process;

    -- Process that verifies the corresponding output
   process
      file inputsFile : text is "test.input"; 
      variable input, expectedOutput : line; 
      variable testCounter : integer := 1;
      variable errorCounter : integer := 0;
      variable expectedOutputString : string(1 to 10000);
      variable testSuccess: boolean;
   begin
      wait for 12 ns; -- wait for reset 
      readline(inputsFile, input); -- skip the first line of advertising
      while not endfile(inputsFile) loop
         readline(inputsFile, input); -- input comment, unused
         readline(inputsFile, input); -- input line, unused
         readline(inputsFile, expectedOutput); -- comment line, unused in this process
         readline(inputsFile, expectedOutput);
         expectedOutputString := expectedOutput.all & (expectedOutput'Length+1 to 10000 => ' ');
         testSuccess := testLine(testCounter, expectedOutputString, expectedOutput'Length, R);
         if not testSuccess then 
               errorCounter := errorCounter + 1; -- incrementing global error counter
         end if;
            testCounter := testCounter + 1; -- incrementing global error counter
         wait for 10 ns;
      end loop;
      report integer'image(errorCounter) & " error(s) encoutered." severity note;
      report "End of simulation after " & integer'image(testCounter-1) & " tests" severity note;
   end process;

end architecture;

