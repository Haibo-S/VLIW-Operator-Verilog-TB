--------------------------------------------------------------------------------
--                          InvA0Table_Freq500_uid8
-- VHDL generated for DummyFPGA @ 500MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 2
-- Target frequency (MHz): 500
-- Input signals: X
-- Output signals: Y
--  approx. input signal timings: X: (c0, 0.000000ns)
--  approx. output signal timings: Y: (c0, 0.550000ns)

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity InvA0Table_Freq500_uid8 is
    port (X : in  std_logic_vector(8 downto 0);
          Y : out  std_logic_vector(9 downto 0)   );
end entity;

architecture arch of InvA0Table_Freq500_uid8 is
signal Y0 :  std_logic_vector(9 downto 0);
   -- timing of Y0: (c0, 0.550000ns)
signal Y1 :  std_logic_vector(9 downto 0);
   -- timing of Y1: (c0, 0.550000ns)
begin
   with X  select  Y0 <= 
      "1000000000" when "000000000",
      "1000000000" when "000000001",
      "0111111111" when "000000010",
      "0111111110" when "000000011",
      "0111111101" when "000000100",
      "0111111100" when "000000101",
      "0111111011" when "000000110",
      "0111111010" when "000000111",
      "0111111001" when "000001000",
      "0111111000" when "000001001",
      "0111110111" when "000001010",
      "0111110110" when "000001011",
      "0111110101" when "000001100",
      "0111110100" when "000001101",
      "0111110011" when "000001110",
      "0111110010" when "000001111",
      "0111110001" when "000010000",
      "0111110000" when "000010001",
      "0111101111" when "000010010",
      "0111101110" when "000010011",
      "0111101101" when "000010100",
      "0111101100" when "000010101",
      "0111101011" when "000010110",
      "0111101010" when "000010111",
      "0111101010" when "000011000",
      "0111101001" when "000011001",
      "0111101000" when "000011010",
      "0111100111" when "000011011",
      "0111100110" when "000011100",
      "0111100101" when "000011101",
      "0111100100" when "000011110",
      "0111100011" when "000011111",
      "0111100010" when "000100000",
      "0111100001" when "000100001",
      "0111100001" when "000100010",
      "0111100000" when "000100011",
      "0111011111" when "000100100",
      "0111011110" when "000100101",
      "0111011101" when "000100110",
      "0111011100" when "000100111",
      "0111011011" when "000101000",
      "0111011011" when "000101001",
      "0111011010" when "000101010",
      "0111011001" when "000101011",
      "0111011000" when "000101100",
      "0111010111" when "000101101",
      "0111010110" when "000101110",
      "0111010101" when "000101111",
      "0111010101" when "000110000",
      "0111010100" when "000110001",
      "0111010011" when "000110010",
      "0111010010" when "000110011",
      "0111010001" when "000110100",
      "0111010000" when "000110101",
      "0111010000" when "000110110",
      "0111001111" when "000110111",
      "0111001110" when "000111000",
      "0111001101" when "000111001",
      "0111001100" when "000111010",
      "0111001100" when "000111011",
      "0111001011" when "000111100",
      "0111001010" when "000111101",
      "0111001001" when "000111110",
      "0111001000" when "000111111",
      "0111001000" when "001000000",
      "0111000111" when "001000001",
      "0111000110" when "001000010",
      "0111000101" when "001000011",
      "0111000100" when "001000100",
      "0111000100" when "001000101",
      "0111000011" when "001000110",
      "0111000010" when "001000111",
      "0111000001" when "001001000",
      "0111000001" when "001001001",
      "0111000000" when "001001010",
      "0110111111" when "001001011",
      "0110111110" when "001001100",
      "0110111110" when "001001101",
      "0110111101" when "001001110",
      "0110111100" when "001001111",
      "0110111011" when "001010000",
      "0110111011" when "001010001",
      "0110111010" when "001010010",
      "0110111001" when "001010011",
      "0110111000" when "001010100",
      "0110111000" when "001010101",
      "0110110111" when "001010110",
      "0110110110" when "001010111",
      "0110110101" when "001011000",
      "0110110101" when "001011001",
      "0110110100" when "001011010",
      "0110110011" when "001011011",
      "0110110011" when "001011100",
      "0110110010" when "001011101",
      "0110110001" when "001011110",
      "0110110000" when "001011111",
      "0110110000" when "001100000",
      "0110101111" when "001100001",
      "0110101110" when "001100010",
      "0110101110" when "001100011",
      "0110101101" when "001100100",
      "0110101100" when "001100101",
      "0110101011" when "001100110",
      "0110101011" when "001100111",
      "0110101010" when "001101000",
      "0110101001" when "001101001",
      "0110101001" when "001101010",
      "0110101000" when "001101011",
      "0110100111" when "001101100",
      "0110100111" when "001101101",
      "0110100110" when "001101110",
      "0110100101" when "001101111",
      "0110100101" when "001110000",
      "0110100100" when "001110001",
      "0110100011" when "001110010",
      "0110100011" when "001110011",
      "0110100010" when "001110100",
      "0110100001" when "001110101",
      "0110100001" when "001110110",
      "0110100000" when "001110111",
      "0110011111" when "001111000",
      "0110011111" when "001111001",
      "0110011110" when "001111010",
      "0110011101" when "001111011",
      "0110011101" when "001111100",
      "0110011100" when "001111101",
      "0110011011" when "001111110",
      "0110011011" when "001111111",
      "0110011010" when "010000000",
      "0110011001" when "010000001",
      "0110011001" when "010000010",
      "0110011000" when "010000011",
      "0110011000" when "010000100",
      "0110010111" when "010000101",
      "0110010110" when "010000110",
      "0110010110" when "010000111",
      "0110010101" when "010001000",
      "0110010100" when "010001001",
      "0110010100" when "010001010",
      "0110010011" when "010001011",
      "0110010011" when "010001100",
      "0110010010" when "010001101",
      "0110010001" when "010001110",
      "0110010001" when "010001111",
      "0110010000" when "010010000",
      "0110010000" when "010010001",
      "0110001111" when "010010010",
      "0110001110" when "010010011",
      "0110001110" when "010010100",
      "0110001101" when "010010101",
      "0110001100" when "010010110",
      "0110001100" when "010010111",
      "0110001011" when "010011000",
      "0110001011" when "010011001",
      "0110001010" when "010011010",
      "0110001010" when "010011011",
      "0110001001" when "010011100",
      "0110001000" when "010011101",
      "0110001000" when "010011110",
      "0110000111" when "010011111",
      "0110000111" when "010100000",
      "0110000110" when "010100001",
      "0110000101" when "010100010",
      "0110000101" when "010100011",
      "0110000100" when "010100100",
      "0110000100" when "010100101",
      "0110000011" when "010100110",
      "0110000011" when "010100111",
      "0110000010" when "010101000",
      "0110000001" when "010101001",
      "0110000001" when "010101010",
      "0110000000" when "010101011",
      "0110000000" when "010101100",
      "0101111111" when "010101101",
      "0101111111" when "010101110",
      "0101111110" when "010101111",
      "0101111110" when "010110000",
      "0101111101" when "010110001",
      "0101111100" when "010110010",
      "0101111100" when "010110011",
      "0101111011" when "010110100",
      "0101111011" when "010110101",
      "0101111010" when "010110110",
      "0101111010" when "010110111",
      "0101111001" when "010111000",
      "0101111001" when "010111001",
      "0101111000" when "010111010",
      "0101111000" when "010111011",
      "0101110111" when "010111100",
      "0101110110" when "010111101",
      "0101110110" when "010111110",
      "0101110101" when "010111111",
      "0101110101" when "011000000",
      "0101110100" when "011000001",
      "0101110100" when "011000010",
      "0101110011" when "011000011",
      "0101110011" when "011000100",
      "0101110010" when "011000101",
      "0101110010" when "011000110",
      "0101110001" when "011000111",
      "0101110001" when "011001000",
      "0101110000" when "011001001",
      "0101110000" when "011001010",
      "0101101111" when "011001011",
      "0101101111" when "011001100",
      "0101101110" when "011001101",
      "0101101110" when "011001110",
      "0101101101" when "011001111",
      "0101101101" when "011010000",
      "0101101100" when "011010001",
      "0101101100" when "011010010",
      "0101101011" when "011010011",
      "0101101011" when "011010100",
      "0101101010" when "011010101",
      "0101101010" when "011010110",
      "0101101001" when "011010111",
      "0101101001" when "011011000",
      "0101101000" when "011011001",
      "0101101000" when "011011010",
      "0101100111" when "011011011",
      "0101100111" when "011011100",
      "0101100110" when "011011101",
      "0101100110" when "011011110",
      "0101100101" when "011011111",
      "0101100101" when "011100000",
      "0101100100" when "011100001",
      "0101100100" when "011100010",
      "0101100011" when "011100011",
      "0101100011" when "011100100",
      "0101100010" when "011100101",
      "0101100010" when "011100110",
      "0101100001" when "011100111",
      "0101100001" when "011101000",
      "0101100000" when "011101001",
      "0101100000" when "011101010",
      "0101011111" when "011101011",
      "0101011111" when "011101100",
      "0101011110" when "011101101",
      "0101011110" when "011101110",
      "0101011110" when "011101111",
      "0101011101" when "011110000",
      "0101011101" when "011110001",
      "0101011100" when "011110010",
      "0101011100" when "011110011",
      "0101011011" when "011110100",
      "0101011011" when "011110101",
      "0101011010" when "011110110",
      "0101011010" when "011110111",
      "0101011001" when "011111000",
      "0101011001" when "011111001",
      "0101011001" when "011111010",
      "0101011000" when "011111011",
      "0101011000" when "011111100",
      "0101010111" when "011111101",
      "0101010111" when "011111110",
      "0101010110" when "011111111",
      "1010101011" when "100000000",
      "1010101010" when "100000001",
      "1010101001" when "100000010",
      "1010101001" when "100000011",
      "1010101000" when "100000100",
      "1010100111" when "100000101",
      "1010100110" when "100000110",
      "1010100101" when "100000111",
      "1010100100" when "100001000",
      "1010100011" when "100001001",
      "1010100010" when "100001010",
      "1010100010" when "100001011",
      "1010100001" when "100001100",
      "1010100000" when "100001101",
      "1010011111" when "100001110",
      "1010011110" when "100001111",
      "1010011101" when "100010000",
      "1010011100" when "100010001",
      "1010011100" when "100010010",
      "1010011011" when "100010011",
      "1010011010" when "100010100",
      "1010011001" when "100010101",
      "1010011000" when "100010110",
      "1010010111" when "100010111",
      "1010010110" when "100011000",
      "1010010110" when "100011001",
      "1010010101" when "100011010",
      "1010010100" when "100011011",
      "1010010011" when "100011100",
      "1010010010" when "100011101",
      "1010010010" when "100011110",
      "1010010001" when "100011111",
      "1010010000" when "100100000",
      "1010001111" when "100100001",
      "1010001110" when "100100010",
      "1010001101" when "100100011",
      "1010001101" when "100100100",
      "1010001100" when "100100101",
      "1010001011" when "100100110",
      "1010001010" when "100100111",
      "1010001001" when "100101000",
      "1010001001" when "100101001",
      "1010001000" when "100101010",
      "1010000111" when "100101011",
      "1010000110" when "100101100",
      "1010000101" when "100101101",
      "1010000101" when "100101110",
      "1010000100" when "100101111",
      "1010000011" when "100110000",
      "1010000010" when "100110001",
      "1010000001" when "100110010",
      "1010000001" when "100110011",
      "1010000000" when "100110100",
      "1001111111" when "100110101",
      "1001111110" when "100110110",
      "1001111110" when "100110111",
      "1001111101" when "100111000",
      "1001111100" when "100111001",
      "1001111011" when "100111010",
      "1001111010" when "100111011",
      "1001111010" when "100111100",
      "1001111001" when "100111101",
      "1001111000" when "100111110",
      "1001110111" when "100111111",
      "1001110111" when "101000000",
      "1001110110" when "101000001",
      "1001110101" when "101000010",
      "1001110100" when "101000011",
      "1001110100" when "101000100",
      "1001110011" when "101000101",
      "1001110010" when "101000110",
      "1001110001" when "101000111",
      "1001110001" when "101001000",
      "1001110000" when "101001001",
      "1001101111" when "101001010",
      "1001101110" when "101001011",
      "1001101110" when "101001100",
      "1001101101" when "101001101",
      "1001101100" when "101001110",
      "1001101011" when "101001111",
      "1001101011" when "101010000",
      "1001101010" when "101010001",
      "1001101001" when "101010010",
      "1001101001" when "101010011",
      "1001101000" when "101010100",
      "1001100111" when "101010101",
      "1001100110" when "101010110",
      "1001100110" when "101010111",
      "1001100101" when "101011000",
      "1001100100" when "101011001",
      "1001100100" when "101011010",
      "1001100011" when "101011011",
      "1001100010" when "101011100",
      "1001100001" when "101011101",
      "1001100001" when "101011110",
      "1001100000" when "101011111",
      "1001011111" when "101100000",
      "1001011111" when "101100001",
      "1001011110" when "101100010",
      "1001011101" when "101100011",
      "1001011101" when "101100100",
      "1001011100" when "101100101",
      "1001011011" when "101100110",
      "1001011010" when "101100111",
      "1001011010" when "101101000",
      "1001011001" when "101101001",
      "1001011000" when "101101010",
      "1001011000" when "101101011",
      "1001010111" when "101101100",
      "1001010110" when "101101101",
      "1001010110" when "101101110",
      "1001010101" when "101101111",
      "1001010100" when "101110000",
      "1001010100" when "101110001",
      "1001010011" when "101110010",
      "1001010010" when "101110011",
      "1001010010" when "101110100",
      "1001010001" when "101110101",
      "1001010000" when "101110110",
      "1001010000" when "101110111",
      "1001001111" when "101111000",
      "1001001110" when "101111001",
      "1001001110" when "101111010",
      "1001001101" when "101111011",
      "1001001100" when "101111100",
      "1001001100" when "101111101",
      "1001001011" when "101111110",
      "1001001010" when "101111111",
      "1001001010" when "110000000",
      "1001001001" when "110000001",
      "1001001000" when "110000010",
      "1001001000" when "110000011",
      "1001000111" when "110000100",
      "1001000110" when "110000101",
      "1001000110" when "110000110",
      "1001000101" when "110000111",
      "1001000100" when "110001000",
      "1001000100" when "110001001",
      "1001000011" when "110001010",
      "1001000011" when "110001011",
      "1001000010" when "110001100",
      "1001000001" when "110001101",
      "1001000001" when "110001110",
      "1001000000" when "110001111",
      "1000111111" when "110010000",
      "1000111111" when "110010001",
      "1000111110" when "110010010",
      "1000111101" when "110010011",
      "1000111101" when "110010100",
      "1000111100" when "110010101",
      "1000111100" when "110010110",
      "1000111011" when "110010111",
      "1000111010" when "110011000",
      "1000111010" when "110011001",
      "1000111001" when "110011010",
      "1000111001" when "110011011",
      "1000111000" when "110011100",
      "1000110111" when "110011101",
      "1000110111" when "110011110",
      "1000110110" when "110011111",
      "1000110101" when "110100000",
      "1000110101" when "110100001",
      "1000110100" when "110100010",
      "1000110100" when "110100011",
      "1000110011" when "110100100",
      "1000110010" when "110100101",
      "1000110010" when "110100110",
      "1000110001" when "110100111",
      "1000110001" when "110101000",
      "1000110000" when "110101001",
      "1000101111" when "110101010",
      "1000101111" when "110101011",
      "1000101110" when "110101100",
      "1000101110" when "110101101",
      "1000101101" when "110101110",
      "1000101100" when "110101111",
      "1000101100" when "110110000",
      "1000101011" when "110110001",
      "1000101011" when "110110010",
      "1000101010" when "110110011",
      "1000101010" when "110110100",
      "1000101001" when "110110101",
      "1000101000" when "110110110",
      "1000101000" when "110110111",
      "1000100111" when "110111000",
      "1000100111" when "110111001",
      "1000100110" when "110111010",
      "1000100101" when "110111011",
      "1000100101" when "110111100",
      "1000100100" when "110111101",
      "1000100100" when "110111110",
      "1000100011" when "110111111",
      "1000100011" when "111000000",
      "1000100010" when "111000001",
      "1000100001" when "111000010",
      "1000100001" when "111000011",
      "1000100000" when "111000100",
      "1000100000" when "111000101",
      "1000011111" when "111000110",
      "1000011111" when "111000111",
      "1000011110" when "111001000",
      "1000011110" when "111001001",
      "1000011101" when "111001010",
      "1000011100" when "111001011",
      "1000011100" when "111001100",
      "1000011011" when "111001101",
      "1000011011" when "111001110",
      "1000011010" when "111001111",
      "1000011010" when "111010000",
      "1000011001" when "111010001",
      "1000011001" when "111010010",
      "1000011000" when "111010011",
      "1000010111" when "111010100",
      "1000010111" when "111010101",
      "1000010110" when "111010110",
      "1000010110" when "111010111",
      "1000010101" when "111011000",
      "1000010101" when "111011001",
      "1000010100" when "111011010",
      "1000010100" when "111011011",
      "1000010011" when "111011100",
      "1000010011" when "111011101",
      "1000010010" when "111011110",
      "1000010010" when "111011111",
      "1000010001" when "111100000",
      "1000010000" when "111100001",
      "1000010000" when "111100010",
      "1000001111" when "111100011",
      "1000001111" when "111100100",
      "1000001110" when "111100101",
      "1000001110" when "111100110",
      "1000001101" when "111100111",
      "1000001101" when "111101000",
      "1000001100" when "111101001",
      "1000001100" when "111101010",
      "1000001011" when "111101011",
      "1000001011" when "111101100",
      "1000001010" when "111101101",
      "1000001010" when "111101110",
      "1000001001" when "111101111",
      "1000001001" when "111110000",
      "1000001000" when "111110001",
      "1000001000" when "111110010",
      "1000000111" when "111110011",
      "1000000111" when "111110100",
      "1000000110" when "111110101",
      "1000000110" when "111110110",
      "1000000101" when "111110111",
      "1000000101" when "111111000",
      "1000000100" when "111111001",
      "1000000100" when "111111010",
      "1000000011" when "111111011",
      "1000000011" when "111111100",
      "1000000010" when "111111101",
      "1000000010" when "111111110",
      "1000000001" when "111111111",
      "----------" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          LogTable1_Freq500_uid22
-- VHDL generated for DummyFPGA @ 500MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 2
-- Target frequency (MHz): 500
-- Input signals: X
-- Output signals: Y
--  approx. input signal timings: X: (c0, 0.000000ns)
--  approx. output signal timings: Y: (c0, 0.550000ns)

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity LogTable1_Freq500_uid22 is
    port (X : in  std_logic_vector(6 downto 0);
          Y : out  std_logic_vector(32 downto 0)   );
end entity;

architecture arch of LogTable1_Freq500_uid22 is
signal Y0 :  std_logic_vector(32 downto 0);
   -- timing of Y0: (c0, 0.550000ns)
signal Y1 :  std_logic_vector(32 downto 0);
   -- timing of Y1: (c0, 0.550000ns)
begin
   with X  select  Y0 <= 
      "000000010000000000000001000000000" when "0000000",
      "000000110000000000000001000000000" when "0000001",
      "000001010000000000001001000000000" when "0000010",
      "000001110000000000011001000000001" when "0000011",
      "000010010000000000110001000000100" when "0000100",
      "000010110000000001010001000001000" when "0000101",
      "000011010000000001111001000001110" when "0000110",
      "000011110000000010101001000010111" when "0000111",
      "000100010000000011100001000100011" when "0001000",
      "000100110000000100100001000110011" when "0001001",
      "000101010000000101101001001001000" when "0001010",
      "000101110000000110111001001100000" when "0001011",
      "000110010000001000010001001111111" when "0001100",
      "000110110000001001110001010100011" when "0001101",
      "000111010000001011011001011001101" when "0001110",
      "000111110000001101001001011111110" when "0001111",
      "001000010000001111000001100110110" when "0010000",
      "001000110000010001000001101110111" when "0010001",
      "001001010000010011001001110111111" when "0010010",
      "001001110000010101011010000010000" when "0010011",
      "001010010000010111110010001101010" when "0010100",
      "001010110000011010010010011001110" when "0010101",
      "001011010000011100111010100111101" when "0010110",
      "001011110000011111101010110110110" when "0010111",
      "001100010000100010100011000111011" when "0011000",
      "001100110000100101100011011001011" when "0011001",
      "001101010000101000101011101101000" when "0011010",
      "001101110000101011111100000010001" when "0011011",
      "001110010000101111010100011000111" when "0011100",
      "001110110000110010110100110001100" when "0011101",
      "001111010000110110011101001011110" when "0011110",
      "001111110000111010001101101000000" when "0011111",
      "010000010000111110000110000110000" when "0100000",
      "010000110001000010000110100110001" when "0100001",
      "010001010001000110001111001000010" when "0100010",
      "010001110001001010011111101100100" when "0100011",
      "010010010001001110111000010010110" when "0100100",
      "010010110001010011011000111011011" when "0100101",
      "010011010001011000000001100110010" when "0100110",
      "010011110001011100110010010011100" when "0100111",
      "010100010001100001101011000011001" when "0101000",
      "010100110001100110101011110101010" when "0101001",
      "010101010001101011110100101010000" when "0101010",
      "010101110001110001000101100001010" when "0101011",
      "010110010001110110011110011011001" when "0101100",
      "010110110001111011111111010111110" when "0101101",
      "010111010010000001101000010111010" when "0101110",
      "010111110010000111011001011001100" when "0101111",
      "011000010010001101010010011110110" when "0110000",
      "011000110010010011010011100111000" when "0110001",
      "011001010010011001011100110010010" when "0110010",
      "011001110010011111101110000000101" when "0110011",
      "011010010010100110000111010010010" when "0110100",
      "011010110010101100101000100111000" when "0110101",
      "011011010010110011010001111111000" when "0110110",
      "011011110010111010000011011010100" when "0110111",
      "011100010011000000111100111001010" when "0111000",
      "011100110011000111111110011011101" when "0111001",
      "011101010011001111001000000001100" when "0111010",
      "011101110011010110011001101011000" when "0111011",
      "011110010011011101110011011000010" when "0111100",
      "011110110011100101010101001001001" when "0111101",
      "011111010011101100111110111101111" when "0111110",
      "011111110011110100110000110110100" when "0111111",
      "100000000011111000101100110100010" when "1000000",
      "100000100100000000101010110010110" when "1000001",
      "100001000100001000110000110101010" when "1000010",
      "100001100100010000111110111011111" when "1000011",
      "100010000100011001010101000110101" when "1000100",
      "100010100100100001110011010101101" when "1000101",
      "100011000100101010011001101000111" when "1000110",
      "100011100100110011001000000000011" when "1000111",
      "100100000100111011111110011100011" when "1001000",
      "100100100101000100111100111100111" when "1001001",
      "100101000101001110000011100001111" when "1001010",
      "100101100101010111010010001011011" when "1001011",
      "100110000101100000101000111001101" when "1001100",
      "100110100101101010000111101100101" when "1001101",
      "100111000101110011101110100100011" when "1001110",
      "100111100101111101011101100001000" when "1001111",
      "101000000110000111010100100010100" when "1010000",
      "101000100110010001010011101001000" when "1010001",
      "101001000110011011011010110100100" when "1010010",
      "101001100110100101101010000101000" when "1010011",
      "101010000110110000000001011010111" when "1010100",
      "101010100110111010100000110101111" when "1010101",
      "101011000111000101001000010110001" when "1010110",
      "101011100111001111110111111011110" when "1010111",
      "101100000111011010101111100110111" when "1011000",
      "101100100111100101101111010111011" when "1011001",
      "101101000111110000110111001101100" when "1011010",
      "101101100111111100000111001001001" when "1011011",
      "101110001000000111011111001010100" when "1011100",
      "101110101000010010111111010001101" when "1011101",
      "101111001000011110100111011110100" when "1011110",
      "101111101000101010010111110001011" when "1011111",
      "110000001000110110010000001010000" when "1100000",
      "110000101001000010010000101000110" when "1100001",
      "110001001001001110011001001101011" when "1100010",
      "110001101001011010101001111000010" when "1100011",
      "110010001001100111000010101001010" when "1100100",
      "110010101001110011100011100000101" when "1100101",
      "110011001010000000001100011110001" when "1100110",
      "110011101010001100111101100010001" when "1100111",
      "110100001010011001110110101100100" when "1101000",
      "110100101010100110110111111101011" when "1101001",
      "110101001010110100000001010100111" when "1101010",
      "110101101011000001010010110010111" when "1101011",
      "110110001011001110101100010111110" when "1101100",
      "110110101011011100001110000011010" when "1101101",
      "110111001011101001110111110101100" when "1101110",
      "110111101011110111101001101110110" when "1101111",
      "111000001100000101100011101111000" when "1110000",
      "111000101100010011100101110110001" when "1110001",
      "111001001100100001110000000100011" when "1110010",
      "111001101100110000000010011001110" when "1110011",
      "111010001100111110011100110110011" when "1110100",
      "111010101101001100111111011010001" when "1110101",
      "111011001101011011101010000101011" when "1110110",
      "111011101101101010011100110111111" when "1110111",
      "111100001101111001010111110001111" when "1111000",
      "111100101110001000011010110011100" when "1111001",
      "111101001110010111100101111100101" when "1111010",
      "111101101110100110111001001101011" when "1111011",
      "111110001110110110010100100101111" when "1111100",
      "111110101111000101111000000110001" when "1111101",
      "111111001111010101100011101110001" when "1111110",
      "111111101111100101010111011110001" when "1111111",
      "---------------------------------" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                 FixRealKCM_Freq500_uid31_T0_Freq500_uid34
-- VHDL generated for DummyFPGA @ 500MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 2
-- Target frequency (MHz): 500
-- Input signals: X
-- Output signals: Y
--  approx. input signal timings: X: (c0, 0.000000ns)
--  approx. output signal timings: Y: (c0, 0.550000ns)

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity FixRealKCM_Freq500_uid31_T0_Freq500_uid34 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(34 downto 0)   );
end entity;

architecture arch of FixRealKCM_Freq500_uid31_T0_Freq500_uid34 is
signal Y0 :  std_logic_vector(34 downto 0);
   -- timing of Y0: (c0, 0.550000ns)
signal Y1 :  std_logic_vector(34 downto 0);
   -- timing of Y1: (c0, 0.550000ns)
begin
   with X  select  Y0 <= 
      "00000000000000000000000000000000000" when "00000",
      "00000101100010111001000010111111110" when "00001",
      "00001011000101110010000101111111100" when "00010",
      "00010000101000101011001000111111010" when "00011",
      "00010110001011100100001011111111000" when "00100",
      "00011011101110011101001110111110110" when "00101",
      "00100001010001010110010001111110100" when "00110",
      "00100110110100001111010100111110010" when "00111",
      "00101100010111001000010111111110000" when "01000",
      "00110001111010000001011010111101110" when "01001",
      "00110111011100111010011101111101100" when "01010",
      "00111100111111110011100000111101010" when "01011",
      "01000010100010101100100011111100111" when "01100",
      "01001000000101100101100110111100101" when "01101",
      "01001101101000011110101001111100011" when "01110",
      "01010011001011010111101100111100001" when "01111",
      "01011000101110010000101111111011111" when "10000",
      "01011110010001001001110010111011101" when "10001",
      "01100011110100000010110101111011011" when "10010",
      "01101001010110111011111000111011001" when "10011",
      "01101110111001110100111011111010111" when "10100",
      "01110100011100101101111110111010101" when "10101",
      "01111001111111100111000001111010011" when "10110",
      "01111111100010100000000100111010001" when "10111",
      "10000101000101011001000111111001111" when "11000",
      "10001010101000010010001010111001101" when "11001",
      "10010000001011001011001101111001011" when "11010",
      "10010101101110000100010000111001001" when "11011",
      "10011011010000111101010011111000111" when "11100",
      "10100000110011110110010110111000101" when "11101",
      "10100110010110101111011001111000011" when "11110",
      "10101011111001101000011100111000001" when "11111",
      "-----------------------------------" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                 FixRealKCM_Freq500_uid31_T1_Freq500_uid37
-- VHDL generated for DummyFPGA @ 500MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 2
-- Target frequency (MHz): 500
-- Input signals: X
-- Output signals: Y
--  approx. input signal timings: X: (c0, 0.000000ns)
--  approx. output signal timings: Y: (c0, 0.550000ns)

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity FixRealKCM_Freq500_uid31_T1_Freq500_uid37 is
    port (X : in  std_logic_vector(2 downto 0);
          Y : out  std_logic_vector(29 downto 0)   );
end entity;

architecture arch of FixRealKCM_Freq500_uid31_T1_Freq500_uid37 is
signal Y0 :  std_logic_vector(29 downto 0);
   -- timing of Y0: (c0, 0.550000ns)
signal Y1 :  std_logic_vector(29 downto 0);
   -- timing of Y1: (c0, 0.550000ns)
begin
   with X  select  Y0 <= 
      "000000000000000000000000000000" when "000",
      "000101100010111001000011000000" when "001",
      "001011000101110010000101111111" when "010",
      "010000101000101011001000111111" when "011",
      "010110001011100100001011111111" when "100",
      "011011101110011101001110111111" when "101",
      "100001010001010110010001111110" when "110",
      "100110110100001111010100111110" when "111",
      "------------------------------" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                            LZOC_23_Freq500_uid4
-- VHDL generated for DummyFPGA @ 500MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007)
--------------------------------------------------------------------------------
-- Pipeline depth: 3 cycles
-- Clock period (ns): 2
-- Target frequency (MHz): 500
-- Input signals: I OZB
-- Output signals: O
--  approx. input signal timings: I: (c0, 0.550000ns)OZB: (c0, 0.000000ns)
--  approx. output signal timings: O: (c3, 0.410000ns)

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity LZOC_23_Freq500_uid4 is
    port (clk : in std_logic;
          I : in  std_logic_vector(22 downto 0);
          OZB : in  std_logic;
          O : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of LZOC_23_Freq500_uid4 is
signal sozb, sozb_d1, sozb_d2 :  std_logic;
   -- timing of sozb: (c0, 0.000000ns)
signal level5, level5_d1 :  std_logic_vector(30 downto 0);
   -- timing of level5: (c0, 0.550000ns)
signal digit4, digit4_d1, digit4_d2 :  std_logic;
   -- timing of digit4: (c0, 1.590000ns)
signal level4, level4_d1 :  std_logic_vector(14 downto 0);
   -- timing of level4: (c1, 0.340000ns)
signal digit3, digit3_d1 :  std_logic;
   -- timing of digit3: (c1, 1.360000ns)
signal level3 :  std_logic_vector(6 downto 0);
   -- timing of level3: (c2, 0.110000ns)
signal digit2 :  std_logic;
   -- timing of digit2: (c2, 1.110000ns)
signal level2, level2_d1 :  std_logic_vector(2 downto 0);
   -- timing of level2: (c2, 1.660000ns)
signal z :  std_logic_vector(2 downto 0);
   -- timing of z: (c3, 0.410000ns)
signal lowBits :  std_logic_vector(1 downto 0);
   -- timing of lowBits: (c3, 0.410000ns)
signal outHighBits, outHighBits_d1 :  std_logic_vector(2 downto 0);
   -- timing of outHighBits: (c2, 1.110000ns)
signal OZB_d1, OZB_d2, OZB_d3 :  std_logic;
   -- timing of OZB: (c0, 0.000000ns)
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            sozb_d1 <=  sozb;
            sozb_d2 <=  sozb_d1;
            level5_d1 <=  level5;
            digit4_d1 <=  digit4;
            digit4_d2 <=  digit4_d1;
            level4_d1 <=  level4;
            digit3_d1 <=  digit3;
            level2_d1 <=  level2;
            outHighBits_d1 <=  outHighBits;
            OZB_d1 <=  OZB;
            OZB_d2 <=  OZB_d1;
            OZB_d3 <=  OZB_d2;
         end if;
      end process;
   sozb <= OZB;
   -- pad input to the next power of two minus 1
   level5 <= I & (7 downto 0 => not sozb);
   -- Main iteration for large inputs
   digit4<= '1' when level5(30 downto 15) = (15 downto 0 => sozb) else '0';
   level4<= level5_d1(14 downto 0) when digit4_d1='1' else level5_d1(30 downto 16);
   digit3<= '1' when level4(14 downto 7) = (7 downto 0 => sozb_d1) else '0';
   level3<= level4_d1(6 downto 0) when digit3_d1='1' else level4_d1(14 downto 8);
   digit2<= '1' when level3(6 downto 3) = (3 downto 0 => sozb_d2) else '0';
   level2<= level3(2 downto 0) when digit2='1' else level3(6 downto 4);
   -- Finish counting with one LUT
   z <= level2_d1 when OZB_d3='0' else (not level2_d1);
   with z  select  lowBits <= 
      "11" when "000",
      "10" when "001",
      "01" when "010",
      "01" when "011",
      "00" when others;
   outHighBits <= digit4_d2 & digit3_d1 & digit2 & "";
   O <= outHighBits_d1 & lowBits ;
end architecture;

--------------------------------------------------------------------------------
--                    LeftShifter12_by_max_12_Freq500_uid6
-- VHDL generated for DummyFPGA @ 500MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca (2008-2011), Florent de Dinechin (2008-2019)
--------------------------------------------------------------------------------
-- Pipeline depth: 4 cycles
-- Clock period (ns): 2
-- Target frequency (MHz): 500
-- Input signals: X S
-- Output signals: R
--  approx. input signal timings: X: (c0, 1.660000ns)S: (c3, 1.460000ns)
--  approx. output signal timings: R: (c4, 1.406154ns)

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity LeftShifter12_by_max_12_Freq500_uid6 is
    port (clk : in std_logic;
          X : in  std_logic_vector(11 downto 0);
          S : in  std_logic_vector(3 downto 0);
          R : out  std_logic_vector(23 downto 0)   );
end entity;

architecture arch of LeftShifter12_by_max_12_Freq500_uid6 is
signal ps, ps_d1 :  std_logic_vector(3 downto 0);
   -- timing of ps: (c3, 1.460000ns)
signal level0, level0_d1, level0_d2, level0_d3 :  std_logic_vector(11 downto 0);
   -- timing of level0: (c0, 1.660000ns)
signal level1, level1_d1 :  std_logic_vector(12 downto 0);
   -- timing of level1: (c3, 1.460000ns)
signal level2 :  std_logic_vector(14 downto 0);
   -- timing of level2: (c4, 0.440769ns)
signal level3 :  std_logic_vector(18 downto 0);
   -- timing of level3: (c4, 0.440769ns)
signal level4 :  std_logic_vector(26 downto 0);
   -- timing of level4: (c4, 1.406154ns)
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            ps_d1 <=  ps;
            level0_d1 <=  level0;
            level0_d2 <=  level0_d1;
            level0_d3 <=  level0_d2;
            level1_d1 <=  level1;
         end if;
      end process;
   ps<= S;
   level0<= X;
   level1<= level0_d3 & (0 downto 0 => '0') when ps(0)= '1' else     (0 downto 0 => '0') & level0_d3;
   level2<= level1_d1 & (1 downto 0 => '0') when ps_d1(1)= '1' else     (1 downto 0 => '0') & level1_d1;
   level3<= level2 & (3 downto 0 => '0') when ps_d1(2)= '1' else     (3 downto 0 => '0') & level2;
   level4<= level3 & (7 downto 0 => '0') when ps_d1(3)= '1' else     (7 downto 0 => '0') & level3;
   R <= level4(23 downto 0);
end architecture;

--------------------------------------------------------------------------------
--                         IntAdder_27_Freq500_uid12
-- VHDL generated for DummyFPGA @ 500MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin (2008-2016)
--------------------------------------------------------------------------------
-- Pipeline depth: 2 cycles
-- Clock period (ns): 2
-- Target frequency (MHz): 500
-- Input signals: X Y Cin
-- Output signals: R
--  approx. input signal timings: X: (c1, 0.640000ns)Y: (c1, 1.190000ns)Cin: (c0, 0.000000ns)
--  approx. output signal timings: R: (c2, 0.660000ns)

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntAdder_27_Freq500_uid12 is
    port (clk : in std_logic;
          X : in  std_logic_vector(26 downto 0);
          Y : in  std_logic_vector(26 downto 0);
          Cin : in  std_logic;
          R : out  std_logic_vector(26 downto 0)   );
end entity;

architecture arch of IntAdder_27_Freq500_uid12 is
signal Cin_1, Cin_1_d1, Cin_1_d2 :  std_logic;
   -- timing of Cin_1: (c0, 0.000000ns)
signal X_1, X_1_d1 :  std_logic_vector(27 downto 0);
   -- timing of X_1: (c1, 0.640000ns)
signal Y_1, Y_1_d1 :  std_logic_vector(27 downto 0);
   -- timing of Y_1: (c1, 1.190000ns)
signal S_1 :  std_logic_vector(27 downto 0);
   -- timing of S_1: (c2, 0.660000ns)
signal R_1 :  std_logic_vector(26 downto 0);
   -- timing of R_1: (c2, 0.660000ns)
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            Cin_1_d1 <=  Cin_1;
            Cin_1_d2 <=  Cin_1_d1;
            X_1_d1 <=  X_1;
            Y_1_d1 <=  Y_1;
         end if;
      end process;
   Cin_1 <= Cin;
   X_1 <= '0' & X(26 downto 0);
   Y_1 <= '0' & Y(26 downto 0);
   S_1 <= X_1_d1 + Y_1_d1 + Cin_1_d2;
   R_1 <= S_1(26 downto 0);
   R <= R_1 ;
end architecture;

--------------------------------------------------------------------------------
--                         IntAdder_27_Freq500_uid15
-- VHDL generated for DummyFPGA @ 500MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin (2008-2016)
--------------------------------------------------------------------------------
-- Pipeline depth: 3 cycles
-- Clock period (ns): 2
-- Target frequency (MHz): 500
-- Input signals: X Y Cin
-- Output signals: R
--  approx. input signal timings: X: (c2, 0.660000ns)Y: (c2, 1.260000ns)Cin: (c0, 0.000000ns)
--  approx. output signal timings: R: (c3, 0.730000ns)

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntAdder_27_Freq500_uid15 is
    port (clk : in std_logic;
          X : in  std_logic_vector(26 downto 0);
          Y : in  std_logic_vector(26 downto 0);
          Cin : in  std_logic;
          R : out  std_logic_vector(26 downto 0)   );
end entity;

architecture arch of IntAdder_27_Freq500_uid15 is
signal Cin_1, Cin_1_d1, Cin_1_d2, Cin_1_d3 :  std_logic;
   -- timing of Cin_1: (c0, 0.000000ns)
signal X_1, X_1_d1 :  std_logic_vector(27 downto 0);
   -- timing of X_1: (c2, 0.660000ns)
signal Y_1, Y_1_d1 :  std_logic_vector(27 downto 0);
   -- timing of Y_1: (c2, 1.260000ns)
signal S_1 :  std_logic_vector(27 downto 0);
   -- timing of S_1: (c3, 0.730000ns)
signal R_1 :  std_logic_vector(26 downto 0);
   -- timing of R_1: (c3, 0.730000ns)
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            Cin_1_d1 <=  Cin_1;
            Cin_1_d2 <=  Cin_1_d1;
            Cin_1_d3 <=  Cin_1_d2;
            X_1_d1 <=  X_1;
            Y_1_d1 <=  Y_1;
         end if;
      end process;
   Cin_1 <= Cin;
   X_1 <= '0' & X(26 downto 0);
   Y_1 <= '0' & Y(26 downto 0);
   S_1 <= X_1_d1 + Y_1_d1 + Cin_1_d3;
   R_1 <= S_1(26 downto 0);
   R <= R_1 ;
end architecture;

--------------------------------------------------------------------------------
--                         IntAdder_27_Freq500_uid18
-- VHDL generated for DummyFPGA @ 500MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin (2008-2016)
--------------------------------------------------------------------------------
-- Pipeline depth: 6 cycles
-- Clock period (ns): 2
-- Target frequency (MHz): 500
-- Input signals: X Y Cin
-- Output signals: R
--  approx. input signal timings: X: (c3, 0.730000ns)Y: (c5, 0.706154ns)Cin: (c0, 0.000000ns)
--  approx. output signal timings: R: (c6, 1.176154ns)

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntAdder_27_Freq500_uid18 is
    port (clk : in std_logic;
          X : in  std_logic_vector(26 downto 0);
          Y : in  std_logic_vector(26 downto 0);
          Cin : in  std_logic;
          R : out  std_logic_vector(26 downto 0)   );
end entity;

architecture arch of IntAdder_27_Freq500_uid18 is
signal Cin_0, Cin_0_d1, Cin_0_d2, Cin_0_d3, Cin_0_d4, Cin_0_d5, Cin_0_d6 :  std_logic;
   -- timing of Cin_0: (c0, 0.000000ns)
signal X_0, X_0_d1, X_0_d2, X_0_d3 :  std_logic_vector(10 downto 0);
   -- timing of X_0: (c3, 0.730000ns)
signal Y_0, Y_0_d1 :  std_logic_vector(10 downto 0);
   -- timing of Y_0: (c5, 0.706154ns)
signal S_0 :  std_logic_vector(10 downto 0);
   -- timing of S_0: (c6, 0.006154ns)
signal R_0 :  std_logic_vector(9 downto 0);
   -- timing of R_0: (c6, 0.006154ns)
signal Cin_1 :  std_logic;
   -- timing of Cin_1: (c6, 0.006154ns)
signal X_1, X_1_d1, X_1_d2, X_1_d3 :  std_logic_vector(17 downto 0);
   -- timing of X_1: (c3, 0.730000ns)
signal Y_1, Y_1_d1 :  std_logic_vector(17 downto 0);
   -- timing of Y_1: (c5, 0.706154ns)
signal S_1 :  std_logic_vector(17 downto 0);
   -- timing of S_1: (c6, 1.176154ns)
signal R_1 :  std_logic_vector(16 downto 0);
   -- timing of R_1: (c6, 1.176154ns)
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            Cin_0_d1 <=  Cin_0;
            Cin_0_d2 <=  Cin_0_d1;
            Cin_0_d3 <=  Cin_0_d2;
            Cin_0_d4 <=  Cin_0_d3;
            Cin_0_d5 <=  Cin_0_d4;
            Cin_0_d6 <=  Cin_0_d5;
            X_0_d1 <=  X_0;
            X_0_d2 <=  X_0_d1;
            X_0_d3 <=  X_0_d2;
            Y_0_d1 <=  Y_0;
            X_1_d1 <=  X_1;
            X_1_d2 <=  X_1_d1;
            X_1_d3 <=  X_1_d2;
            Y_1_d1 <=  Y_1;
         end if;
      end process;
   Cin_0 <= Cin;
   X_0 <= '0' & X(9 downto 0);
   Y_0 <= '0' & Y(9 downto 0);
   S_0 <= X_0_d3 + Y_0_d1 + Cin_0_d6;
   R_0 <= S_0(9 downto 0);
   Cin_1 <= S_0(10);
   X_1 <= '0' & X(26 downto 10);
   Y_1 <= '0' & Y(26 downto 10);
   S_1 <= X_1_d3 + Y_1_d1 + Cin_1;
   R_1 <= S_1(16 downto 0);
   R <= R_1 & R_0 ;
end architecture;

--------------------------------------------------------------------------------
--                          LogTable0_Freq500_uid20
-- VHDL generated for DummyFPGA @ 500MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- Pipeline depth: 2 cycles
-- Clock period (ns): 2
-- Target frequency (MHz): 500
-- Input signals: X
-- Output signals: Y
--  approx. input signal timings: X: (c0, 0.000000ns)
--  approx. output signal timings: Y: (c2, 0.415625ns)

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity LogTable0_Freq500_uid20 is
    port (clk : in std_logic;
          X : in  std_logic_vector(8 downto 0);
          Y : out  std_logic_vector(39 downto 0)   );
end entity;

architecture arch of LogTable0_Freq500_uid20 is
signal Y0, Y0_d1 :  std_logic_vector(39 downto 0);
   -- timing of Y0: (c1, 0.200000ns)
signal Y1 :  std_logic_vector(39 downto 0);
   -- timing of Y1: (c2, 0.415625ns)
signal X_d1 :  std_logic_vector(8 downto 0);
   -- timing of X: (c0, 0.000000ns)
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            Y0_d1 <=  Y0;
            X_d1 <=  X;
         end if;
      end process;
   with X_d1  select  Y0 <= 
      "1111111111111100000000000000000000000000" when "000000000",
      "1111111111111100000000000000000000000000" when "000000001",
      "0000000001111100001000000000101010101111" when "000000010",
      "0000000011111100100000000101010110010110" when "000000011",
      "0000000101111101001000010010000101000110" when "000000100",
      "0000000111111110000000101010111010110001" when "000000101",
      "0000001001111111001001010011111100101101" when "000000110",
      "0000001100000000100010010001010001110001" when "000000111",
      "0000001110000010001011100111000010011001" when "000001000",
      "0000010000000100000101011001011000100101" when "000001001",
      "0000010010000110001111101100011111111011" when "000001010",
      "0000010100001000101010100100100101100110" when "000001011",
      "0000010110001011010110000101111000011010" when "000001100",
      "0000011000001110010010010100101000110010" when "000001101",
      "0000011010010001011111010101001000110001" when "000001110",
      "0000011100010100111101001011101100000101" when "000001111",
      "0000011110011000101011111100101000000101" when "000010000",
      "0000100000011100101011101100010011110100" when "000010001",
      "0000100010100000111100011111001000000000" when "000010010",
      "0000100100100101011110011001011111000111" when "000010011",
      "0000100110101010010001011111110101010001" when "000010100",
      "0000101000101111010101110110101000010111" when "000010101",
      "0000101010110100101011100010011000000010" when "000010110",
      "0000101100111010010010100111100101101010" when "000010111",
      "0000101100111010010010100111100101101010" when "000011000",
      "0000101111000000001011001010110100011011" when "000011001",
      "0000110001000110010101010000101001010000" when "000011010",
      "0000110011001100110000111101101010111010" when "000011011",
      "0000110101010011011110010110100001111110" when "000011100",
      "0000110111011010011101011111111000110100" when "000011101",
      "0000111001100001101110011110011011101111" when "000011110",
      "0000111011101001010001010110111000110100" when "000011111",
      "0000111101110001000110001110000000000011" when "000100000",
      "0000111111111001001101001000100011010110" when "000100001",
      "0000111111111001001101001000100011010110" when "000100010",
      "0001000010000001100110001011010110011110" when "000100011",
      "0001000100001010010001011011001111001011" when "000100100",
      "0001000110010011001110111101000101000110" when "000100101",
      "0001001000011100011110110101110001111000" when "000100110",
      "0001001010100110000001001010010001000111" when "000100111",
      "0001001100101111110101111111100000011000" when "000101000",
      "0001001100101111110101111111100000011000" when "000101001",
      "0001001110111001111101011010011111010010" when "000101010",
      "0001010001000100010111100000001111011100" when "000101011",
      "0001010011001111000100010101110100100000" when "000101100",
      "0001010101011010000100000000010100001110" when "000101101",
      "0001010111100101010110100100110110011000" when "000101110",
      "0001011001110000111100001000100100110110" when "000101111",
      "0001011001110000111100001000100100110110" when "000110000",
      "0001011011111100110100110000101011101011" when "000110001",
      "0001011110001001000000100010011000111110" when "000110010",
      "0001100000010101011111100010111101000001" when "000110011",
      "0001100010100010010001110111101010010010" when "000110100",
      "0001100100101111010111100101110101011001" when "000110101",
      "0001100100101111010111100101110101011001" when "000110110",
      "0001100110111100110000110010110101001101" when "000110111",
      "0001101001001010011101100100000010110010" when "000111000",
      "0001101011011000011101111110111001011011" when "000111001",
      "0001101101100110110010001000110110101101" when "000111010",
      "0001101101100110110010001000110110101101" when "000111011",
      "0001101111110101011010000111011010100000" when "000111100",
      "0001110010000100010110000000000110111100" when "000111101",
      "0001110100010011100101111000100000100010" when "000111110",
      "0001110110100011001001110110001110000100" when "000111111",
      "0001110110100011001001110110001110000100" when "001000000",
      "0001111000110011000001111110111000110000" when "001000001",
      "0001111011000011001110011000001100001010" when "001000010",
      "0001111101010011101111000111110110010000" when "001000011",
      "0001111111100100100100010011100111011100" when "001000100",
      "0001111111100100100100010011100111011100" when "001000101",
      "0010000001110101101110000001010010100100" when "001000110",
      "0010000100000111001100010110101100111100" when "001000111",
      "0010000110011000111111011001101110011010" when "001001000",
      "0010000110011000111111011001101110011010" when "001001001",
      "0010001000101011000111010000010001010000" when "001001010",
      "0010001010111101100100000000010010010110" when "001001011",
      "0010001101010000010101101111110001001000" when "001001100",
      "0010001101010000010101101111110001001000" when "001001101",
      "0010001111100011011100100100101111100101" when "001001110",
      "0010010001110110111000100101010010010100" when "001001111",
      "0010010100001010101001110111100000100011" when "001010000",
      "0010010100001010101001110111100000100011" when "001010001",
      "0010010110011110110000100001100100001101" when "001010010",
      "0010011000110011001100101001101001110100" when "001010011",
      "0010011011000111111110010110000000101011" when "001010100",
      "0010011011000111111110010110000000101011" when "001010101",
      "0010011101011101000101101100111010110000" when "001010110",
      "0010011111110010100010110100101100110010" when "001010111",
      "0010100010001000010101110011101110010100" when "001011000",
      "0010100010001000010101110011101110010100" when "001011001",
      "0010100100011110011110110000011001101000" when "001011010",
      "0010100110110100111101110001001011111000" when "001011011",
      "0010100110110100111101110001001011111000" when "001011100",
      "0010101001001011110010111100100101000100" when "001011101",
      "0010101011100010111110011001001000000011" when "001011110",
      "0010101101111010100000001101011010101000" when "001011111",
      "0010101101111010100000001101011010101000" when "001100000",
      "0010110000010010011000100000000101100001" when "001100001",
      "0010110010101010100111010111110100011000" when "001100010",
      "0010110010101010100111010111110100011000" when "001100011",
      "0010110101000011001100111011010101111000" when "001100100",
      "0010110111011100001001010001011011101011" when "001100101",
      "0010111001110101011100100000111010100000" when "001100110",
      "0010111001110101011100100000111010100000" when "001100111",
      "0010111100001111000110110000101010001000" when "001101000",
      "0010111110101001001000000111100101011111" when "001101001",
      "0010111110101001001000000111100101011111" when "001101010",
      "0011000001000011100000101100101010100011" when "001101011",
      "0011000011011110010000100110111010100010" when "001101100",
      "0011000011011110010000100110111010100010" when "001101101",
      "0011000101111001010111111101011001110010" when "001101110",
      "0011001000010100110110110111001111111010" when "001101111",
      "0011001000010100110110110111001111111010" when "001110000",
      "0011001010110000101101011011100111101110" when "001110001",
      "0011001101001100111011110001101111010111" when "001110010",
      "0011001101001100111011110001101111010111" when "001110011",
      "0011001111101001100010000000111000010001" when "001110100",
      "0011010010000110100000010000010111001101" when "001110101",
      "0011010010000110100000010000010111001101" when "001110110",
      "0011010100100011110110100111100100010110" when "001110111",
      "0011010111000001100101001101111011001110" when "001111000",
      "0011010111000001100101001101111011001110" when "001111001",
      "0011011001011111101100001010111010111000" when "001111010",
      "0011011011111110001011100110000101110000" when "001111011",
      "0011011011111110001011100110000101110000" when "001111100",
      "0011011110011101000011100111000001111000" when "001111101",
      "0011100000111100010100010101011000110000" when "001111110",
      "0011100000111100010100010101011000110000" when "001111111",
      "0011100011011011111101111000110111100000" when "010000000",
      "0011100101111100000000011001001110110110" when "010000001",
      "0011100101111100000000011001001110110110" when "010000010",
      "0011101000011100011011111110010011001011" when "010000011",
      "0011101000011100011011111110010011001011" when "010000100",
      "0011101010111101010000101111111100100000" when "010000101",
      "0011101101011110011110110110000110101001" when "010000110",
      "0011101101011110011110110110000110101001" when "010000111",
      "0011110000000000000110011000110001000111" when "010001000",
      "0011110010100010000111011111111111001110" when "010001001",
      "0011110010100010000111011111111111001110" when "010001010",
      "0011110101000100100010010011111000001001" when "010001011",
      "0011110101000100100010010011111000001001" when "010001100",
      "0011110111100111010110111100100110111010" when "010001101",
      "0011111010001010100101100010011010011100" when "010001110",
      "0011111010001010100101100010011010011100" when "010001111",
      "0011111100101110001110001101100101101000" when "010010000",
      "0011111100101110001110001101100101101000" when "010010001",
      "0011111111010010010001000110011111010100" when "010010010",
      "0100000001110110101110010101100010011011" when "010010011",
      "0100000001110110101110010101100010011011" when "010010100",
      "0100000100011011100110000011001101111010" when "010010101",
      "0100000111000000111000011000000100110110" when "010010110",
      "0100000111000000111000011000000100110110" when "010010111",
      "0100001001100110100101011100101110011011" when "010011000",
      "0100001001100110100101011100101110011011" when "010011001",
      "0100001100001100101101011001110110000110" when "010011010",
      "0100001100001100101101011001110110000110" when "010011011",
      "0100001110110011010000011000001011011110" when "010011100",
      "0100010001011010001110100000100010100000" when "010011101",
      "0100010001011010001110100000100010100000" when "010011110",
      "0100010100000001100111111011110011011010" when "010011111",
      "0100010100000001100111111011110011011010" when "010100000",
      "0100010110101001011100110010111010110100" when "010100001",
      "0100011001010001101101001110111001101111" when "010100010",
      "0100011001010001101101001110111001101111" when "010100011",
      "0100011011111010011001011000110101101010" when "010100100",
      "0100011011111010011001011000110101101010" when "010100101",
      "0100011110100011100001011001111000100010" when "010100110",
      "0100011110100011100001011001111000100010" when "010100111",
      "0100100001001101000101011011010000111011" when "010101000",
      "0100100011110111000101100110010001111011" when "010101001",
      "0100100011110111000101100110010001111011" when "010101010",
      "0100100110100001100010000100010011010100" when "010101011",
      "0100100110100001100010000100010011010100" when "010101100",
      "0100101001001100011010111110110001100010" when "010101101",
      "0100101001001100011010111110110001100010" when "010101110",
      "0100101011110111110000011111001101110010" when "010101111",
      "0100101011110111110000011111001101110010" when "010110000",
      "0100101110100011100010101111001110000100" when "010110001",
      "0100110001001111110001111000011101001110" when "010110010",
      "0100110001001111110001111000011101001110" when "010110011",
      "0100110011111100011110000100101010111011" when "010110100",
      "0100110011111100011110000100101010111011" when "010110101",
      "0100110110101001100111011101101011111000" when "010110110",
      "0100110110101001100111011101101011111000" when "010110111",
      "0100111001010111001110001101011001101111" when "010111000",
      "0100111001010111001110001101011001101111" when "010111001",
      "0100111100000101010010011101110011001101" when "010111010",
      "0100111100000101010010011101110011001101" when "010111011",
      "0100111110110011110100011000111100000110" when "010111100",
      "0101000001100010110100001000111101011000" when "010111101",
      "0101000001100010110100001000111101011000" when "010111110",
      "0101000100010010010001111000000101001110" when "010111111",
      "0101000100010010010001111000000101001110" when "011000000",
      "0101000111000010001101110000100111000111" when "011000001",
      "0101000111000010001101110000100111000111" when "011000010",
      "0101001001110010100111111100111011110011" when "011000011",
      "0101001001110010100111111100111011110011" when "011000100",
      "0101001100100011100000100111100001011100" when "011000101",
      "0101001100100011100000100111100001011100" when "011000110",
      "0101001111010100110111111010111011101010" when "011000111",
      "0101001111010100110111111010111011101010" when "011001000",
      "0101010010000110101110000001110011100010" when "011001001",
      "0101010010000110101110000001110011100010" when "011001010",
      "0101010100111001000011000110110111110000" when "011001011",
      "0101010100111001000011000110110111110000" when "011001100",
      "0101010111101011110111010100111100100100" when "011001101",
      "0101010111101011110111010100111100100100" when "011001110",
      "0101011010011111001010110110111011111100" when "011001111",
      "0101011010011111001010110110111011111100" when "011010000",
      "0101011101010010111101110111110101100110" when "011010001",
      "0101011101010010111101110111110101100110" when "011010010",
      "0101100000000111010000100010101111000010" when "011010011",
      "0101100000000111010000100010101111000010" when "011010100",
      "0101100010111100000011000010110011101010" when "011010101",
      "0101100010111100000011000010110011101010" when "011010110",
      "0101100101110001010101100011010100110100" when "011010111",
      "0101100101110001010101100011010100110100" when "011011000",
      "0101101000100111001000001111101001110010" when "011011001",
      "0101101000100111001000001111101001110010" when "011011010",
      "0101101011011101011011010011001111111110" when "011011011",
      "0101101011011101011011010011001111111110" when "011011100",
      "0101101110010100001110111001101010111100" when "011011101",
      "0101101110010100001110111001101010111100" when "011011110",
      "0101110001001011100011001110100100011010" when "011011111",
      "0101110001001011100011001110100100011010" when "011100000",
      "0101110100000011011000011101101100011010" when "011100001",
      "0101110100000011011000011101101100011010" when "011100010",
      "0101110110111011101110110010111001010010" when "011100011",
      "0101110110111011101110110010111001010010" when "011100100",
      "0101111001110100100110011010000111110100" when "011100101",
      "0101111001110100100110011010000111110100" when "011100110",
      "0101111100101101111111011111011011010010" when "011100111",
      "0101111100101101111111011111011011010010" when "011101000",
      "0101111111100111111010001110111101100000" when "011101001",
      "0101111111100111111010001110111101100000" when "011101010",
      "0110000010100010010110110100111110111110" when "011101011",
      "0110000010100010010110110100111110111110" when "011101100",
      "0110000101011101010101011101110110110111" when "011101101",
      "0110000101011101010101011101110110110111" when "011101110",
      "0110000101011101010101011101110110110111" when "011101111",
      "0110001000011000110110010110000011001010" when "011110000",
      "0110001000011000110110010110000011001010" when "011110001",
      "0110001011010100111001101010001000101100" when "011110010",
      "0110001011010100111001101010001000101100" when "011110011",
      "0110001110010001011111100110110011010010" when "011110100",
      "0110001110010001011111100110110011010010" when "011110101",
      "0110010001001110101000011000110101110000" when "011110110",
      "0110010001001110101000011000110101110000" when "011110111",
      "0110010100001100010100001101001010000001" when "011111000",
      "0110010100001100010100001101001010000001" when "011111001",
      "0110010100001100010100001101001010000001" when "011111010",
      "0110010111001010100011010000110001001110" when "011111011",
      "0110010111001010100011010000110001001110" when "011111100",
      "0110011010001001010101110000110011110000" when "011111101",
      "0110011010001001010101110000110011110000" when "011111110",
      "0110011101001000101011111010100001011000" when "011111111",
      "1011011000110110011110011011101100000010" when "100000000",
      "1011011010010110011111111011110010000010" when "100000001",
      "1011011011110110101010011101000000001100" when "100000010",
      "1011011011110110101010011101000000001100" when "100000011",
      "1011011101010110111110000001000011000010" when "100000100",
      "1011011110110111011010101001100111101000" when "100000101",
      "1011100000011000000000011000011011011110" when "100000110",
      "1011100001111000101111001111001100100100" when "100000111",
      "1011100011011001100111001111101001011010" when "100001000",
      "1011100100111010101000011011100000111110" when "100001001",
      "1011100110011011110010110100100010110000" when "100001010",
      "1011100110011011110010110100100010110000" when "100001011",
      "1011100111111101000110011100011110101100" when "100001100",
      "1011101001011110100011010101000101010010" when "100001101",
      "1011101011000000001001100000000111011110" when "100001110",
      "1011101100100001111000111111010110110010" when "100001111",
      "1011101110000011110001110100100101001010" when "100010000",
      "1011101111100101110100000001100101000111" when "100010001",
      "1011101111100101110100000001100101000111" when "100010010",
      "1011110001000111111111101000001001101010" when "100010011",
      "1011110010101010010100101010000110010101" when "100010100",
      "1011110100001100110011001001001111001100" when "100010101",
      "1011110101101111011011000111011000110010" when "100010110",
      "1011110111010010001100100110011000001110" when "100010111",
      "1011111000110101000111101000000011001010" when "100011000",
      "1011111000110101000111101000000011001010" when "100011001",
      "1011111010011000001100001110001111110000" when "100011010",
      "1011111011111011011010011010110100101100" when "100011011",
      "1011111101011110110010001111101001010000" when "100011100",
      "1011111111000010010011101110100101001010" when "100011101",
      "1011111111000010010011101110100101001010" when "100011110",
      "1100000000100101111110111001100000110100" when "100011111",
      "1100000010001001110011110010010101000100" when "100100000",
      "1100000011101101110010011010111011010101" when "100100001",
      "1100000101010001111010110101001101101001" when "100100010",
      "1100000110110110001101000011000110100010" when "100100011",
      "1100000110110110001101000011000110100010" when "100100100",
      "1100001000011010101001000110100001000111" when "100100101",
      "1100001001111111001111000001011001000101" when "100100110",
      "1100001011100011111110110101101010101011" when "100100111",
      "1100001101001000111000100101010010101111" when "100101000",
      "1100001101001000111000100101010010101111" when "100101001",
      "1100001110101101111100010010001110101010" when "100101010",
      "1100010000010011001001111110011100011100" when "100101011",
      "1100010001111000100001101011111010101000" when "100101100",
      "1100010011011110000011011100101000011010" when "100101101",
      "1100010011011110000011011100101000011010" when "100101110",
      "1100010101000011101111010010100101100000" when "100101111",
      "1100010110101001100101001111110010010010" when "100110000",
      "1100011000001111100101010110001111101100" when "100110001",
      "1100011001110101101111100111111111010001" when "100110010",
      "1100011001110101101111100111111111010001" when "100110011",
      "1100011011011100000100000111000011001011" when "100110100",
      "1100011101000010100010110101011110001010" when "100110101",
      "1100011110101001001011110101010011101000" when "100110110",
      "1100011110101001001011110101010011101000" when "100110111",
      "1100100000001111111111001000100111100100" when "100111000",
      "1100100001110110111100110001011110100101" when "100111001",
      "1100100011011110000100110001111101111100" when "100111010",
      "1100100101000101010111001100001011100000" when "100111011",
      "1100100101000101010111001100001011100000" when "100111100",
      "1100100110101100110100000010001101110100" when "100111101",
      "1100101000010100011011010110001011111110" when "100111110",
      "1100101001111100001101001010001101110100" when "100111111",
      "1100101001111100001101001010001101110100" when "101000000",
      "1100101011100100001001100000011011110000" when "101000001",
      "1100101101001100010000011010111110111000" when "101000010",
      "1100101110110100100001111100000000111010" when "101000011",
      "1100101110110100100001111100000000111010" when "101000100",
      "1100110000011100111110000101101100010011" when "101000101",
      "1100110010000101100100111010001100000100" when "101000110",
      "1100110011101110010110011011101011111101" when "101000111",
      "1100110011101110010110011011101011111101" when "101001000",
      "1100110101010111010010101100011000010111" when "101001001",
      "1100110111000000011001101110011110011000" when "101001010",
      "1100111000101001101011100100001011101111" when "101001011",
      "1100111000101001101011100100001011101111" when "101001100",
      "1100111010010011001000001111101110111001" when "101001101",
      "1100111011111100101111110011010110111110" when "101001110",
      "1100111101100110100010010001010011110011" when "101001111",
      "1100111101100110100010010001010011110011" when "101010000",
      "1100111111010000011111101011110101111001" when "101010001",
      "1101000000111010101000000101001110011110" when "101010010",
      "1101000000111010101000000101001110011110" when "101010011",
      "1101000010100100111011011111101111011110" when "101010100",
      "1101000100001111011001111101101011100010" when "101010101",
      "1101000101111010000011100001010110000000" when "101010110",
      "1101000101111010000011100001010110000000" when "101010111",
      "1101000111100100111000001101000010111101" when "101011000",
      "1101001001001111111000000011000111001100" when "101011001",
      "1101001001001111111000000011000111001100" when "101011010",
      "1101001010111011000011000101111000010001" when "101011011",
      "1101001100100110011001010111101100011011" when "101011100",
      "1101001110010001111010111010111010101011" when "101011101",
      "1101001110010001111010111010111010101011" when "101011110",
      "1101001111111101100111110001111010110001" when "101011111",
      "1101010001101001011111111111000101001101" when "101100000",
      "1101010001101001011111111111000101001101" when "101100001",
      "1101010011010101100011100100110011010000" when "101100010",
      "1101010101000001110010100101011110111010" when "101100011",
      "1101010101000001110010100101011110111010" when "101100100",
      "1101010110101110001101000011100010111100" when "101100101",
      "1101011000011010110011000001011010111100" when "101100110",
      "1101011010000111100100100001100011001011" when "101100111",
      "1101011010000111100100100001100011001011" when "101101000",
      "1101011011110100100001100110011000110010" when "101101001",
      "1101011101100001101010010010011001101001" when "101101010",
      "1101011101100001101010010010011001101001" when "101101011",
      "1101011111001110111110101000000100011011" when "101101100",
      "1101100000111100011110101001111000100110" when "101101101",
      "1101100000111100011110101001111000100110" when "101101110",
      "1101100010101010001010011010010110011101" when "101101111",
      "1101100100011000000001111011111111000011" when "101110000",
      "1101100100011000000001111011111111000011" when "101110001",
      "1101100110000110000101010001010100010010" when "101110010",
      "1101100111110100010100011100111000110111" when "101110011",
      "1101100111110100010100011100111000110111" when "101110100",
      "1101101001100010101111100001010000010100" when "101110101",
      "1101101011010001010110100000111111000000" when "101110110",
      "1101101011010001010110100000111111000000" when "101110111",
      "1101101101000000001001011110101010000111" when "101111000",
      "1101101110101111001000011100110111101011" when "101111001",
      "1101101110101111001000011100110111101011" when "101111010",
      "1101110000011110010011011110001110100100" when "101111011",
      "1101110010001101101010100101010110100001" when "101111100",
      "1101110010001101101010100101010110100001" when "101111101",
      "1101110011111101001101110100111000000111" when "101111110",
      "1101110101101100111101001111011100110010" when "101111111",
      "1101110101101100111101001111011100110010" when "110000000",
      "1101110111011100111000110111101110110110" when "110000001",
      "1101111001001101000000110000011001011111" when "110000010",
      "1101111001001101000000110000011001011111" when "110000011",
      "1101111010111101010100111100001000110010" when "110000100",
      "1101111100101101110101011101101001101011" when "110000101",
      "1101111100101101110101011101101001101011" when "110000110",
      "1101111110011110100010010111101010000010" when "110000111",
      "1110000000001111011011101100111000100100" when "110001000",
      "1110000000001111011011101100111000100100" when "110001001",
      "1110000010000000100001100000000100111100" when "110001010",
      "1110000010000000100001100000000100111100" when "110001011",
      "1110000011110001110011110011111111101111" when "110001100",
      "1110000101100011010010101011011010011001" when "110001101",
      "1110000101100011010010101011011010011001" when "110001110",
      "1110000111010100111110001001000111010101" when "110001111",
      "1110001001000110110110001111111001111000" when "110010000",
      "1110001001000110110110001111111001111000" when "110010001",
      "1110001010111000111011000010100110010011" when "110010010",
      "1110001100101011001100100100000001110100" when "110010011",
      "1110001100101011001100100100000001110100" when "110010100",
      "1110001110011101101010110111000010100100" when "110010101",
      "1110001110011101101010110111000010100100" when "110010110",
      "1110010000010000010101111110011111101100" when "110010111",
      "1110010010000011001101111101010001001111" when "110011000",
      "1110010010000011001101111101010001001111" when "110011001",
      "1110010011110110010010110110010000010010" when "110011010",
      "1110010011110110010010110110010000010010" when "110011011",
      "1110010101101001100100101100010110110101" when "110011100",
      "1110010111011101000011100010011111111010" when "110011101",
      "1110010111011101000011100010011111111010" when "110011110",
      "1110011001010000101111011011100111100000" when "110011111",
      "1110011011000100101000011010101010100111" when "110100000",
      "1110011011000100101000011010101010100111" when "110100001",
      "1110011100111000101110100010100111001110" when "110100010",
      "1110011100111000101110100010100111001110" when "110100011",
      "1110011110101101000001110110011100011000" when "110100100",
      "1110100000100001100010011001001010000101" when "110100101",
      "1110100000100001100010011001001010000101" when "110100110",
      "1110100010010110010000001101110001011001" when "110100111",
      "1110100010010110010000001101110001011001" when "110101000",
      "1110100100001011001011010111010100011011" when "110101001",
      "1110100110000000010011111000110110010001" when "110101010",
      "1110100110000000010011111000110110010001" when "110101011",
      "1110100111110101101001110101011011001001" when "110101100",
      "1110100111110101101001110101011011001001" when "110101101",
      "1110101001101011001101010000001000010000" when "110101110",
      "1110101011100000111110001100000011111010" when "110101111",
      "1110101011100000111110001100000011111010" when "110110000",
      "1110101101010110111100101100010101011110" when "110110001",
      "1110101101010110111100101100010101011110" when "110110010",
      "1110101111001101001000110100000101011010" when "110110011",
      "1110101111001101001000110100000101011010" when "110110100",
      "1110110001000011100010100110011101001110" when "110110101",
      "1110110010111010001010000110100111100100" when "110110110",
      "1110110010111010001010000110100111100100" when "110110111",
      "1110110100110000111111010111110000001010" when "110111000",
      "1110110100110000111111010111110000001010" when "110111001",
      "1110110110101000000010011101000011110110" when "110111010",
      "1110111000011111010011011001110000100101" when "110111011",
      "1110111000011111010011011001110000100101" when "110111100",
      "1110111010010110110010010001000101011100" when "110111101",
      "1110111010010110110010010001000101011100" when "110111110",
      "1110111100001110011111000110010010101011" when "110111111",
      "1110111100001110011111000110010010101011" when "111000000",
      "1110111110000110011001111100101001100111" when "111000001",
      "1110111111111110100010110111011100110010" when "111000010",
      "1110111111111110100010110111011100110010" when "111000011",
      "1111000001110110111001111001111111110111" when "111000100",
      "1111000001110110111001111001111111110111" when "111000101",
      "1111000011101111011111000111100111101100" when "111000110",
      "1111000011101111011111000111100111101100" when "111000111",
      "1111000101101000010010100011101010010010" when "111001000",
      "1111000101101000010010100011101010010010" when "111001001",
      "1111000111100001010100010001011110110111" when "111001010",
      "1111001001011010100100010100011101110011" when "111001011",
      "1111001001011010100100010100011101110011" when "111001100",
      "1111001011010100000010110000000000101110" when "111001101",
      "1111001011010100000010110000000000101110" when "111001110",
      "1111001101001101101111100111100010011100" when "111001111",
      "1111001101001101101111100111100010011100" when "111010000",
      "1111001111000111101010111110011110111110" when "111010001",
      "1111001111000111101010111110011110111110" when "111010010",
      "1111010001000001110100111000010011100111" when "111010011",
      "1111010010111100001101011000011110110110" when "111010100",
      "1111010010111100001101011000011110110110" when "111010101",
      "1111010100110110110100100010100000011100" when "111010110",
      "1111010100110110110100100010100000011100" when "111010111",
      "1111010110110001101010011001111001011001" when "111011000",
      "1111010110110001101010011001111001011001" when "111011001",
      "1111011000101100101111000010001100000001" when "111011010",
      "1111011000101100101111000010001100000001" when "111011011",
      "1111011010101000000010011110111011110110" when "111011100",
      "1111011010101000000010011110111011110110" when "111011101",
      "1111011100100011100100110011101101101110" when "111011110",
      "1111011100100011100100110011101101101110" when "111011111",
      "1111011110011111010110000100000111110011" when "111100000",
      "1111100000011011010110010011110001100010" when "111100001",
      "1111100000011011010110010011110001100010" when "111100010",
      "1111100010010111100101100110010011101011" when "111100011",
      "1111100010010111100101100110010011101011" when "111100100",
      "1111100100010100000011111111011000010100" when "111100101",
      "1111100100010100000011111111011000010100" when "111100110",
      "1111100110010000110001100010101010111001" when "111100111",
      "1111100110010000110001100010101010111001" when "111101000",
      "1111101000001101101110010011111000001011" when "111101001",
      "1111101000001101101110010011111000001011" when "111101010",
      "1111101010001010111010010110101110010010" when "111101011",
      "1111101010001010111010010110101110010010" when "111101100",
      "1111101100001000010101101110111100101110" when "111101101",
      "1111101100001000010101101110111100101110" when "111101110",
      "1111101110000110000000100000010100011000" when "111101111",
      "1111101110000110000000100000010100011000" when "111110000",
      "1111110000000011111010101110100111100000" when "111110001",
      "1111110000000011111010101110100111100000" when "111110010",
      "1111110010000010000100011101101001110001" when "111110011",
      "1111110010000010000100011101101001110001" when "111110100",
      "1111110100000000011101110001010000010000" when "111110101",
      "1111110100000000011101110001010000010000" when "111110110",
      "1111110101111111000110101101010001011011" when "111110111",
      "1111110101111111000110101101010001011011" when "111111000",
      "1111110111111101111111010101100101001111" when "111111001",
      "1111110111111101111111010101100101001111" when "111111010",
      "1111111001111101000111101110000101000010" when "111111011",
      "1111111001111101000111101110000101000010" when "111111100",
      "1111111011111100011111111010101011101010" when "111111101",
      "1111111011111100011111111010101011101010" when "111111110",
      "1111111101111100000111111111010101011001" when "111111111",
      "----------------------------------------" when others;
   Y1 <= Y0_d1; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                         IntAdder_40_Freq500_uid26
-- VHDL generated for DummyFPGA @ 500MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin (2008-2016)
--------------------------------------------------------------------------------
-- Pipeline depth: 3 cycles
-- Clock period (ns): 2
-- Target frequency (MHz): 500
-- Input signals: X Y Cin
-- Output signals: R
--  approx. input signal timings: X: (c2, 0.415625ns)Y: (c1, 1.190000ns)Cin: (c0, 0.000000ns)
--  approx. output signal timings: R: (c3, 1.015625ns)

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntAdder_40_Freq500_uid26 is
    port (clk : in std_logic;
          X : in  std_logic_vector(39 downto 0);
          Y : in  std_logic_vector(39 downto 0);
          Cin : in  std_logic;
          R : out  std_logic_vector(39 downto 0)   );
end entity;

architecture arch of IntAdder_40_Freq500_uid26 is
signal Cin_0, Cin_0_d1, Cin_0_d2, Cin_0_d3 :  std_logic;
   -- timing of Cin_0: (c0, 0.000000ns)
signal X_0, X_0_d1 :  std_logic_vector(39 downto 0);
   -- timing of X_0: (c2, 0.415625ns)
signal Y_0, Y_0_d1, Y_0_d2 :  std_logic_vector(39 downto 0);
   -- timing of Y_0: (c1, 1.190000ns)
signal S_0 :  std_logic_vector(39 downto 0);
   -- timing of S_0: (c3, 0.005625ns)
signal R_0 :  std_logic_vector(38 downto 0);
   -- timing of R_0: (c3, 0.005625ns)
signal Cin_1 :  std_logic;
   -- timing of Cin_1: (c3, 0.005625ns)
signal X_1, X_1_d1 :  std_logic_vector(1 downto 0);
   -- timing of X_1: (c2, 0.415625ns)
signal Y_1, Y_1_d1, Y_1_d2 :  std_logic_vector(1 downto 0);
   -- timing of Y_1: (c1, 1.190000ns)
signal S_1 :  std_logic_vector(1 downto 0);
   -- timing of S_1: (c3, 1.015625ns)
signal R_1 :  std_logic_vector(0 downto 0);
   -- timing of R_1: (c3, 1.015625ns)
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            Cin_0_d1 <=  Cin_0;
            Cin_0_d2 <=  Cin_0_d1;
            Cin_0_d3 <=  Cin_0_d2;
            X_0_d1 <=  X_0;
            Y_0_d1 <=  Y_0;
            Y_0_d2 <=  Y_0_d1;
            X_1_d1 <=  X_1;
            Y_1_d1 <=  Y_1;
            Y_1_d2 <=  Y_1_d1;
         end if;
      end process;
   Cin_0 <= Cin;
   X_0 <= '0' & X(38 downto 0);
   Y_0 <= '0' & Y(38 downto 0);
   S_0 <= X_0_d1 + Y_0_d2 + Cin_0_d3;
   R_0 <= S_0(38 downto 0);
   Cin_1 <= S_0(39);
   X_1 <= '0' & X(39 downto 39);
   Y_1 <= '0' & Y(39 downto 39);
   S_1 <= X_1_d1 + Y_1_d2 + Cin_1;
   R_1 <= S_1(0 downto 0);
   R <= R_1 & R_0 ;
end architecture;

--------------------------------------------------------------------------------
--                         IntAdder_40_Freq500_uid29
-- VHDL generated for DummyFPGA @ 500MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin (2008-2016)
--------------------------------------------------------------------------------
-- Pipeline depth: 7 cycles
-- Clock period (ns): 2
-- Target frequency (MHz): 500
-- Input signals: X Y Cin
-- Output signals: R
--  approx. input signal timings: X: (c3, 1.015625ns)Y: (c6, 1.176154ns)Cin: (c0, 0.000000ns)
--  approx. output signal timings: R: (c7, 0.776154ns)

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntAdder_40_Freq500_uid29 is
    port (clk : in std_logic;
          X : in  std_logic_vector(39 downto 0);
          Y : in  std_logic_vector(39 downto 0);
          Cin : in  std_logic;
          R : out  std_logic_vector(39 downto 0)   );
end entity;

architecture arch of IntAdder_40_Freq500_uid29 is
signal Cin_1, Cin_1_d1, Cin_1_d2, Cin_1_d3, Cin_1_d4, Cin_1_d5, Cin_1_d6, Cin_1_d7 :  std_logic;
   -- timing of Cin_1: (c0, 0.000000ns)
signal X_1, X_1_d1, X_1_d2, X_1_d3, X_1_d4 :  std_logic_vector(40 downto 0);
   -- timing of X_1: (c3, 1.015625ns)
signal Y_1, Y_1_d1 :  std_logic_vector(40 downto 0);
   -- timing of Y_1: (c6, 1.176154ns)
signal S_1 :  std_logic_vector(40 downto 0);
   -- timing of S_1: (c7, 0.776154ns)
signal R_1 :  std_logic_vector(39 downto 0);
   -- timing of R_1: (c7, 0.776154ns)
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            Cin_1_d1 <=  Cin_1;
            Cin_1_d2 <=  Cin_1_d1;
            Cin_1_d3 <=  Cin_1_d2;
            Cin_1_d4 <=  Cin_1_d3;
            Cin_1_d5 <=  Cin_1_d4;
            Cin_1_d6 <=  Cin_1_d5;
            Cin_1_d7 <=  Cin_1_d6;
            X_1_d1 <=  X_1;
            X_1_d2 <=  X_1_d1;
            X_1_d3 <=  X_1_d2;
            X_1_d4 <=  X_1_d3;
            Y_1_d1 <=  Y_1;
         end if;
      end process;
   Cin_1 <= Cin;
   X_1 <= '0' & X(39 downto 0);
   Y_1 <= '0' & Y(39 downto 0);
   S_1 <= X_1_d4 + Y_1_d1 + Cin_1_d7;
   R_1 <= S_1(39 downto 0);
   R <= R_1 ;
end architecture;

--------------------------------------------------------------------------------
--                         IntAdder_35_Freq500_uid41
-- VHDL generated for DummyFPGA @ 500MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin (2008-2016)
--------------------------------------------------------------------------------
-- Pipeline depth: 1 cycles
-- Clock period (ns): 2
-- Target frequency (MHz): 500
-- Input signals: X Y Cin
-- Output signals: R
--  approx. input signal timings: X: (c1, 0.370000ns)Y: (c1, 0.370000ns)Cin: (c0, 0.000000ns)
--  approx. output signal timings: R: (c1, 1.710000ns)

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntAdder_35_Freq500_uid41 is
    port (clk : in std_logic;
          X : in  std_logic_vector(34 downto 0);
          Y : in  std_logic_vector(34 downto 0);
          Cin : in  std_logic;
          R : out  std_logic_vector(34 downto 0)   );
end entity;

architecture arch of IntAdder_35_Freq500_uid41 is
signal Rtmp :  std_logic_vector(34 downto 0);
   -- timing of Rtmp: (c1, 1.710000ns)
signal Cin_d1 :  std_logic;
   -- timing of Cin: (c0, 0.000000ns)
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            Cin_d1 <=  Cin;
         end if;
      end process;
   Rtmp <= X + Y + Cin_d1;
   R <= Rtmp;
end architecture;

--------------------------------------------------------------------------------
--                          FixRealKCM_Freq500_uid31
-- VHDL generated for DummyFPGA @ 500MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin (2007-2016)
--------------------------------------------------------------------------------
-- Pipeline depth: 1 cycles
-- Clock period (ns): 2
-- Target frequency (MHz): 500
-- Input signals: X
-- Output signals: R
--  approx. input signal timings: X: (c0, 1.620000ns)
--  approx. output signal timings: R: (c1, 1.710000ns)

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity FixRealKCM_Freq500_uid31 is
    port (clk : in std_logic;
          X : in  std_logic_vector(7 downto 0);
          R : out  std_logic_vector(34 downto 0)   );
end entity;

architecture arch of FixRealKCM_Freq500_uid31 is
   component FixRealKCM_Freq500_uid31_T0_Freq500_uid34 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(34 downto 0)   );
   end component;

   component FixRealKCM_Freq500_uid31_T1_Freq500_uid37 is
      port ( X : in  std_logic_vector(2 downto 0);
             Y : out  std_logic_vector(29 downto 0)   );
   end component;

   component IntAdder_35_Freq500_uid41 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(34 downto 0);
             Y : in  std_logic_vector(34 downto 0);
             Cin : in  std_logic;
             R : out  std_logic_vector(34 downto 0)   );
   end component;

signal FixRealKCM_Freq500_uid31_A0 :  std_logic_vector(4 downto 0);
   -- timing of FixRealKCM_Freq500_uid31_A0: (c0, 1.620000ns)
signal FixRealKCM_Freq500_uid31_T0 :  std_logic_vector(34 downto 0);
   -- timing of FixRealKCM_Freq500_uid31_T0: (c1, 0.370000ns)
signal FixRealKCM_Freq500_uid31_T0_copy35, FixRealKCM_Freq500_uid31_T0_copy35_d1 :  std_logic_vector(34 downto 0);
   -- timing of FixRealKCM_Freq500_uid31_T0_copy35: (c0, 1.620000ns)
signal bh32_w0_0 :  std_logic;
   -- timing of bh32_w0_0: (c1, 0.370000ns)
signal bh32_w1_0 :  std_logic;
   -- timing of bh32_w1_0: (c1, 0.370000ns)
signal bh32_w2_0 :  std_logic;
   -- timing of bh32_w2_0: (c1, 0.370000ns)
signal bh32_w3_0 :  std_logic;
   -- timing of bh32_w3_0: (c1, 0.370000ns)
signal bh32_w4_0 :  std_logic;
   -- timing of bh32_w4_0: (c1, 0.370000ns)
signal bh32_w5_0 :  std_logic;
   -- timing of bh32_w5_0: (c1, 0.370000ns)
signal bh32_w6_0 :  std_logic;
   -- timing of bh32_w6_0: (c1, 0.370000ns)
signal bh32_w7_0 :  std_logic;
   -- timing of bh32_w7_0: (c1, 0.370000ns)
signal bh32_w8_0 :  std_logic;
   -- timing of bh32_w8_0: (c1, 0.370000ns)
signal bh32_w9_0 :  std_logic;
   -- timing of bh32_w9_0: (c1, 0.370000ns)
signal bh32_w10_0 :  std_logic;
   -- timing of bh32_w10_0: (c1, 0.370000ns)
signal bh32_w11_0 :  std_logic;
   -- timing of bh32_w11_0: (c1, 0.370000ns)
signal bh32_w12_0 :  std_logic;
   -- timing of bh32_w12_0: (c1, 0.370000ns)
signal bh32_w13_0 :  std_logic;
   -- timing of bh32_w13_0: (c1, 0.370000ns)
signal bh32_w14_0 :  std_logic;
   -- timing of bh32_w14_0: (c1, 0.370000ns)
signal bh32_w15_0 :  std_logic;
   -- timing of bh32_w15_0: (c1, 0.370000ns)
signal bh32_w16_0 :  std_logic;
   -- timing of bh32_w16_0: (c1, 0.370000ns)
signal bh32_w17_0 :  std_logic;
   -- timing of bh32_w17_0: (c1, 0.370000ns)
signal bh32_w18_0 :  std_logic;
   -- timing of bh32_w18_0: (c1, 0.370000ns)
signal bh32_w19_0 :  std_logic;
   -- timing of bh32_w19_0: (c1, 0.370000ns)
signal bh32_w20_0 :  std_logic;
   -- timing of bh32_w20_0: (c1, 0.370000ns)
signal bh32_w21_0 :  std_logic;
   -- timing of bh32_w21_0: (c1, 0.370000ns)
signal bh32_w22_0 :  std_logic;
   -- timing of bh32_w22_0: (c1, 0.370000ns)
signal bh32_w23_0 :  std_logic;
   -- timing of bh32_w23_0: (c1, 0.370000ns)
signal bh32_w24_0 :  std_logic;
   -- timing of bh32_w24_0: (c1, 0.370000ns)
signal bh32_w25_0 :  std_logic;
   -- timing of bh32_w25_0: (c1, 0.370000ns)
signal bh32_w26_0 :  std_logic;
   -- timing of bh32_w26_0: (c1, 0.370000ns)
signal bh32_w27_0 :  std_logic;
   -- timing of bh32_w27_0: (c1, 0.370000ns)
signal bh32_w28_0 :  std_logic;
   -- timing of bh32_w28_0: (c1, 0.370000ns)
signal bh32_w29_0 :  std_logic;
   -- timing of bh32_w29_0: (c1, 0.370000ns)
signal bh32_w30_0 :  std_logic;
   -- timing of bh32_w30_0: (c1, 0.370000ns)
signal bh32_w31_0 :  std_logic;
   -- timing of bh32_w31_0: (c1, 0.370000ns)
signal bh32_w32_0 :  std_logic;
   -- timing of bh32_w32_0: (c1, 0.370000ns)
signal bh32_w33_0 :  std_logic;
   -- timing of bh32_w33_0: (c1, 0.370000ns)
signal bh32_w34_0 :  std_logic;
   -- timing of bh32_w34_0: (c1, 0.370000ns)
signal FixRealKCM_Freq500_uid31_A1 :  std_logic_vector(2 downto 0);
   -- timing of FixRealKCM_Freq500_uid31_A1: (c0, 1.620000ns)
signal FixRealKCM_Freq500_uid31_T1 :  std_logic_vector(29 downto 0);
   -- timing of FixRealKCM_Freq500_uid31_T1: (c1, 0.370000ns)
signal FixRealKCM_Freq500_uid31_T1_copy38, FixRealKCM_Freq500_uid31_T1_copy38_d1 :  std_logic_vector(29 downto 0);
   -- timing of FixRealKCM_Freq500_uid31_T1_copy38: (c0, 1.620000ns)
signal bh32_w0_1 :  std_logic;
   -- timing of bh32_w0_1: (c1, 0.370000ns)
signal bh32_w1_1 :  std_logic;
   -- timing of bh32_w1_1: (c1, 0.370000ns)
signal bh32_w2_1 :  std_logic;
   -- timing of bh32_w2_1: (c1, 0.370000ns)
signal bh32_w3_1 :  std_logic;
   -- timing of bh32_w3_1: (c1, 0.370000ns)
signal bh32_w4_1 :  std_logic;
   -- timing of bh32_w4_1: (c1, 0.370000ns)
signal bh32_w5_1 :  std_logic;
   -- timing of bh32_w5_1: (c1, 0.370000ns)
signal bh32_w6_1 :  std_logic;
   -- timing of bh32_w6_1: (c1, 0.370000ns)
signal bh32_w7_1 :  std_logic;
   -- timing of bh32_w7_1: (c1, 0.370000ns)
signal bh32_w8_1 :  std_logic;
   -- timing of bh32_w8_1: (c1, 0.370000ns)
signal bh32_w9_1 :  std_logic;
   -- timing of bh32_w9_1: (c1, 0.370000ns)
signal bh32_w10_1 :  std_logic;
   -- timing of bh32_w10_1: (c1, 0.370000ns)
signal bh32_w11_1 :  std_logic;
   -- timing of bh32_w11_1: (c1, 0.370000ns)
signal bh32_w12_1 :  std_logic;
   -- timing of bh32_w12_1: (c1, 0.370000ns)
signal bh32_w13_1 :  std_logic;
   -- timing of bh32_w13_1: (c1, 0.370000ns)
signal bh32_w14_1 :  std_logic;
   -- timing of bh32_w14_1: (c1, 0.370000ns)
signal bh32_w15_1 :  std_logic;
   -- timing of bh32_w15_1: (c1, 0.370000ns)
signal bh32_w16_1 :  std_logic;
   -- timing of bh32_w16_1: (c1, 0.370000ns)
signal bh32_w17_1 :  std_logic;
   -- timing of bh32_w17_1: (c1, 0.370000ns)
signal bh32_w18_1 :  std_logic;
   -- timing of bh32_w18_1: (c1, 0.370000ns)
signal bh32_w19_1 :  std_logic;
   -- timing of bh32_w19_1: (c1, 0.370000ns)
signal bh32_w20_1 :  std_logic;
   -- timing of bh32_w20_1: (c1, 0.370000ns)
signal bh32_w21_1 :  std_logic;
   -- timing of bh32_w21_1: (c1, 0.370000ns)
signal bh32_w22_1 :  std_logic;
   -- timing of bh32_w22_1: (c1, 0.370000ns)
signal bh32_w23_1 :  std_logic;
   -- timing of bh32_w23_1: (c1, 0.370000ns)
signal bh32_w24_1 :  std_logic;
   -- timing of bh32_w24_1: (c1, 0.370000ns)
signal bh32_w25_1 :  std_logic;
   -- timing of bh32_w25_1: (c1, 0.370000ns)
signal bh32_w26_1 :  std_logic;
   -- timing of bh32_w26_1: (c1, 0.370000ns)
signal bh32_w27_1 :  std_logic;
   -- timing of bh32_w27_1: (c1, 0.370000ns)
signal bh32_w28_1 :  std_logic;
   -- timing of bh32_w28_1: (c1, 0.370000ns)
signal bh32_w29_1 :  std_logic;
   -- timing of bh32_w29_1: (c1, 0.370000ns)
signal bitheapFinalAdd_bh32_In0 :  std_logic_vector(34 downto 0);
   -- timing of bitheapFinalAdd_bh32_In0: (c1, 0.370000ns)
signal bitheapFinalAdd_bh32_In1 :  std_logic_vector(34 downto 0);
   -- timing of bitheapFinalAdd_bh32_In1: (c1, 0.370000ns)
signal bitheapFinalAdd_bh32_Cin :  std_logic;
   -- timing of bitheapFinalAdd_bh32_Cin: (c0, 0.000000ns)
signal bitheapFinalAdd_bh32_Out :  std_logic_vector(34 downto 0);
   -- timing of bitheapFinalAdd_bh32_Out: (c1, 1.710000ns)
signal bitheapResult_bh32 :  std_logic_vector(34 downto 0);
   -- timing of bitheapResult_bh32: (c1, 1.710000ns)
signal OutRes :  std_logic_vector(34 downto 0);
   -- timing of OutRes: (c1, 1.710000ns)
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            FixRealKCM_Freq500_uid31_T0_copy35_d1 <=  FixRealKCM_Freq500_uid31_T0_copy35;
            FixRealKCM_Freq500_uid31_T1_copy38_d1 <=  FixRealKCM_Freq500_uid31_T1_copy38;
         end if;
      end process;
-- This operator multiplies by log(2)
   FixRealKCM_Freq500_uid31_A0 <= X(7 downto 3);-- input address  m=7  l=3
   FixRealKCM_Freq500_uid31_Table0: FixRealKCM_Freq500_uid31_T0_Freq500_uid34
      port map ( X => FixRealKCM_Freq500_uid31_A0,
                 Y => FixRealKCM_Freq500_uid31_T0_copy35);
   FixRealKCM_Freq500_uid31_T0 <= FixRealKCM_Freq500_uid31_T0_copy35_d1; -- output copy to hold a pipeline register if needed
   bh32_w0_0 <= FixRealKCM_Freq500_uid31_T0(0);
   bh32_w1_0 <= FixRealKCM_Freq500_uid31_T0(1);
   bh32_w2_0 <= FixRealKCM_Freq500_uid31_T0(2);
   bh32_w3_0 <= FixRealKCM_Freq500_uid31_T0(3);
   bh32_w4_0 <= FixRealKCM_Freq500_uid31_T0(4);
   bh32_w5_0 <= FixRealKCM_Freq500_uid31_T0(5);
   bh32_w6_0 <= FixRealKCM_Freq500_uid31_T0(6);
   bh32_w7_0 <= FixRealKCM_Freq500_uid31_T0(7);
   bh32_w8_0 <= FixRealKCM_Freq500_uid31_T0(8);
   bh32_w9_0 <= FixRealKCM_Freq500_uid31_T0(9);
   bh32_w10_0 <= FixRealKCM_Freq500_uid31_T0(10);
   bh32_w11_0 <= FixRealKCM_Freq500_uid31_T0(11);
   bh32_w12_0 <= FixRealKCM_Freq500_uid31_T0(12);
   bh32_w13_0 <= FixRealKCM_Freq500_uid31_T0(13);
   bh32_w14_0 <= FixRealKCM_Freq500_uid31_T0(14);
   bh32_w15_0 <= FixRealKCM_Freq500_uid31_T0(15);
   bh32_w16_0 <= FixRealKCM_Freq500_uid31_T0(16);
   bh32_w17_0 <= FixRealKCM_Freq500_uid31_T0(17);
   bh32_w18_0 <= FixRealKCM_Freq500_uid31_T0(18);
   bh32_w19_0 <= FixRealKCM_Freq500_uid31_T0(19);
   bh32_w20_0 <= FixRealKCM_Freq500_uid31_T0(20);
   bh32_w21_0 <= FixRealKCM_Freq500_uid31_T0(21);
   bh32_w22_0 <= FixRealKCM_Freq500_uid31_T0(22);
   bh32_w23_0 <= FixRealKCM_Freq500_uid31_T0(23);
   bh32_w24_0 <= FixRealKCM_Freq500_uid31_T0(24);
   bh32_w25_0 <= FixRealKCM_Freq500_uid31_T0(25);
   bh32_w26_0 <= FixRealKCM_Freq500_uid31_T0(26);
   bh32_w27_0 <= FixRealKCM_Freq500_uid31_T0(27);
   bh32_w28_0 <= FixRealKCM_Freq500_uid31_T0(28);
   bh32_w29_0 <= FixRealKCM_Freq500_uid31_T0(29);
   bh32_w30_0 <= FixRealKCM_Freq500_uid31_T0(30);
   bh32_w31_0 <= FixRealKCM_Freq500_uid31_T0(31);
   bh32_w32_0 <= FixRealKCM_Freq500_uid31_T0(32);
   bh32_w33_0 <= FixRealKCM_Freq500_uid31_T0(33);
   bh32_w34_0 <= FixRealKCM_Freq500_uid31_T0(34);
   FixRealKCM_Freq500_uid31_A1 <= X(2 downto 0);-- input address  m=2  l=0
   FixRealKCM_Freq500_uid31_Table1: FixRealKCM_Freq500_uid31_T1_Freq500_uid37
      port map ( X => FixRealKCM_Freq500_uid31_A1,
                 Y => FixRealKCM_Freq500_uid31_T1_copy38);
   FixRealKCM_Freq500_uid31_T1 <= FixRealKCM_Freq500_uid31_T1_copy38_d1; -- output copy to hold a pipeline register if needed
   bh32_w0_1 <= FixRealKCM_Freq500_uid31_T1(0);
   bh32_w1_1 <= FixRealKCM_Freq500_uid31_T1(1);
   bh32_w2_1 <= FixRealKCM_Freq500_uid31_T1(2);
   bh32_w3_1 <= FixRealKCM_Freq500_uid31_T1(3);
   bh32_w4_1 <= FixRealKCM_Freq500_uid31_T1(4);
   bh32_w5_1 <= FixRealKCM_Freq500_uid31_T1(5);
   bh32_w6_1 <= FixRealKCM_Freq500_uid31_T1(6);
   bh32_w7_1 <= FixRealKCM_Freq500_uid31_T1(7);
   bh32_w8_1 <= FixRealKCM_Freq500_uid31_T1(8);
   bh32_w9_1 <= FixRealKCM_Freq500_uid31_T1(9);
   bh32_w10_1 <= FixRealKCM_Freq500_uid31_T1(10);
   bh32_w11_1 <= FixRealKCM_Freq500_uid31_T1(11);
   bh32_w12_1 <= FixRealKCM_Freq500_uid31_T1(12);
   bh32_w13_1 <= FixRealKCM_Freq500_uid31_T1(13);
   bh32_w14_1 <= FixRealKCM_Freq500_uid31_T1(14);
   bh32_w15_1 <= FixRealKCM_Freq500_uid31_T1(15);
   bh32_w16_1 <= FixRealKCM_Freq500_uid31_T1(16);
   bh32_w17_1 <= FixRealKCM_Freq500_uid31_T1(17);
   bh32_w18_1 <= FixRealKCM_Freq500_uid31_T1(18);
   bh32_w19_1 <= FixRealKCM_Freq500_uid31_T1(19);
   bh32_w20_1 <= FixRealKCM_Freq500_uid31_T1(20);
   bh32_w21_1 <= FixRealKCM_Freq500_uid31_T1(21);
   bh32_w22_1 <= FixRealKCM_Freq500_uid31_T1(22);
   bh32_w23_1 <= FixRealKCM_Freq500_uid31_T1(23);
   bh32_w24_1 <= FixRealKCM_Freq500_uid31_T1(24);
   bh32_w25_1 <= FixRealKCM_Freq500_uid31_T1(25);
   bh32_w26_1 <= FixRealKCM_Freq500_uid31_T1(26);
   bh32_w27_1 <= FixRealKCM_Freq500_uid31_T1(27);
   bh32_w28_1 <= FixRealKCM_Freq500_uid31_T1(28);
   bh32_w29_1 <= FixRealKCM_Freq500_uid31_T1(29);

   -- Adding the constant bits 
      -- All the constant bits are zero, nothing to add


   bitheapFinalAdd_bh32_In0 <= "" & bh32_w34_0 & bh32_w33_0 & bh32_w32_0 & bh32_w31_0 & bh32_w30_0 & bh32_w29_1 & bh32_w28_1 & bh32_w27_1 & bh32_w26_1 & bh32_w25_1 & bh32_w24_1 & bh32_w23_1 & bh32_w22_1 & bh32_w21_1 & bh32_w20_1 & bh32_w19_1 & bh32_w18_1 & bh32_w17_1 & bh32_w16_1 & bh32_w15_1 & bh32_w14_1 & bh32_w13_1 & bh32_w12_1 & bh32_w11_1 & bh32_w10_1 & bh32_w9_1 & bh32_w8_1 & bh32_w7_1 & bh32_w6_1 & bh32_w5_1 & bh32_w4_1 & bh32_w3_1 & bh32_w2_1 & bh32_w1_1 & bh32_w0_1;
   bitheapFinalAdd_bh32_In1 <= "0" & "0" & "0" & "0" & "0" & bh32_w29_0 & bh32_w28_0 & bh32_w27_0 & bh32_w26_0 & bh32_w25_0 & bh32_w24_0 & bh32_w23_0 & bh32_w22_0 & bh32_w21_0 & bh32_w20_0 & bh32_w19_0 & bh32_w18_0 & bh32_w17_0 & bh32_w16_0 & bh32_w15_0 & bh32_w14_0 & bh32_w13_0 & bh32_w12_0 & bh32_w11_0 & bh32_w10_0 & bh32_w9_0 & bh32_w8_0 & bh32_w7_0 & bh32_w6_0 & bh32_w5_0 & bh32_w4_0 & bh32_w3_0 & bh32_w2_0 & bh32_w1_0 & bh32_w0_0;
   bitheapFinalAdd_bh32_Cin <= '0';

   bitheapFinalAdd_bh32: IntAdder_35_Freq500_uid41
      port map ( clk  => clk,
                 Cin => bitheapFinalAdd_bh32_Cin,
                 X => bitheapFinalAdd_bh32_In0,
                 Y => bitheapFinalAdd_bh32_In1,
                 R => bitheapFinalAdd_bh32_Out);
   bitheapResult_bh32 <= bitheapFinalAdd_bh32_Out(34 downto 0);
   OutRes <= bitheapResult_bh32(34 downto 0);
   R <= OutRes(34 downto 0);
end architecture;

--------------------------------------------------------------------------------
--                         IntAdder_48_Freq500_uid43
-- VHDL generated for DummyFPGA @ 500MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin (2008-2016)
--------------------------------------------------------------------------------
-- Pipeline depth: 8 cycles
-- Clock period (ns): 2
-- Target frequency (MHz): 500
-- Input signals: X Y Cin
-- Output signals: R
--  approx. input signal timings: X: (c1, 1.710000ns)Y: (c7, 0.776154ns)Cin: (c0, 0.550000ns)
--  approx. output signal timings: R: (c8, 1.456154ns)

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntAdder_48_Freq500_uid43 is
    port (clk : in std_logic;
          X : in  std_logic_vector(47 downto 0);
          Y : in  std_logic_vector(47 downto 0);
          Cin : in  std_logic;
          R : out  std_logic_vector(47 downto 0)   );
end entity;

architecture arch of IntAdder_48_Freq500_uid43 is
signal Cin_0, Cin_0_d1, Cin_0_d2, Cin_0_d3, Cin_0_d4, Cin_0_d5, Cin_0_d6, Cin_0_d7, Cin_0_d8 :  std_logic;
   -- timing of Cin_0: (c0, 0.550000ns)
signal X_0, X_0_d1, X_0_d2, X_0_d3, X_0_d4, X_0_d5, X_0_d6, X_0_d7 :  std_logic_vector(3 downto 0);
   -- timing of X_0: (c1, 1.710000ns)
signal Y_0, Y_0_d1 :  std_logic_vector(3 downto 0);
   -- timing of Y_0: (c7, 0.776154ns)
signal S_0 :  std_logic_vector(3 downto 0);
   -- timing of S_0: (c8, 0.006154ns)
signal R_0 :  std_logic_vector(2 downto 0);
   -- timing of R_0: (c8, 0.006154ns)
signal Cin_1 :  std_logic;
   -- timing of Cin_1: (c8, 0.006154ns)
signal X_1, X_1_d1, X_1_d2, X_1_d3, X_1_d4, X_1_d5, X_1_d6, X_1_d7 :  std_logic_vector(45 downto 0);
   -- timing of X_1: (c1, 1.710000ns)
signal Y_1, Y_1_d1 :  std_logic_vector(45 downto 0);
   -- timing of Y_1: (c7, 0.776154ns)
signal S_1 :  std_logic_vector(45 downto 0);
   -- timing of S_1: (c8, 1.456154ns)
signal R_1 :  std_logic_vector(44 downto 0);
   -- timing of R_1: (c8, 1.456154ns)
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            Cin_0_d1 <=  Cin_0;
            Cin_0_d2 <=  Cin_0_d1;
            Cin_0_d3 <=  Cin_0_d2;
            Cin_0_d4 <=  Cin_0_d3;
            Cin_0_d5 <=  Cin_0_d4;
            Cin_0_d6 <=  Cin_0_d5;
            Cin_0_d7 <=  Cin_0_d6;
            Cin_0_d8 <=  Cin_0_d7;
            X_0_d1 <=  X_0;
            X_0_d2 <=  X_0_d1;
            X_0_d3 <=  X_0_d2;
            X_0_d4 <=  X_0_d3;
            X_0_d5 <=  X_0_d4;
            X_0_d6 <=  X_0_d5;
            X_0_d7 <=  X_0_d6;
            Y_0_d1 <=  Y_0;
            X_1_d1 <=  X_1;
            X_1_d2 <=  X_1_d1;
            X_1_d3 <=  X_1_d2;
            X_1_d4 <=  X_1_d3;
            X_1_d5 <=  X_1_d4;
            X_1_d6 <=  X_1_d5;
            X_1_d7 <=  X_1_d6;
            Y_1_d1 <=  Y_1;
         end if;
      end process;
   Cin_0 <= Cin;
   X_0 <= '0' & X(2 downto 0);
   Y_0 <= '0' & Y(2 downto 0);
   S_0 <= X_0_d7 + Y_0_d1 + Cin_0_d8;
   R_0 <= S_0(2 downto 0);
   Cin_1 <= S_0(3);
   X_1 <= '0' & X(47 downto 3);
   Y_1 <= '0' & Y(47 downto 3);
   S_1 <= X_1_d7 + Y_1_d1 + Cin_1;
   R_1 <= S_1(44 downto 0);
   R <= R_1 & R_0 ;
end architecture;

--------------------------------------------------------------------------------
--                    Normalizer_Z_48_40_19_Freq500_uid45
-- VHDL generated for DummyFPGA @ 500MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, (2007-2020)
--------------------------------------------------------------------------------
-- Pipeline depth: 3 cycles
-- Clock period (ns): 2
-- Target frequency (MHz): 500
-- Input signals: X
-- Output signals: Count R
--  approx. input signal timings: X: (c8, 1.456154ns)
--  approx. output signal timings: Count: (c11, 1.096154ns)R: (c11, 1.646154ns)

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity Normalizer_Z_48_40_19_Freq500_uid45 is
    port (clk : in std_logic;
          X : in  std_logic_vector(47 downto 0);
          Count : out  std_logic_vector(4 downto 0);
          R : out  std_logic_vector(39 downto 0)   );
end entity;

architecture arch of Normalizer_Z_48_40_19_Freq500_uid45 is
signal level5, level5_d1 :  std_logic_vector(47 downto 0);
   -- timing of level5: (c8, 1.456154ns)
signal count4, count4_d1, count4_d2 :  std_logic;
   -- timing of count4: (c9, 0.246154ns)
signal level4, level4_d1 :  std_logic_vector(47 downto 0);
   -- timing of level4: (c9, 0.796154ns)
signal count3, count3_d1, count3_d2 :  std_logic;
   -- timing of count3: (c9, 1.366154ns)
signal level3 :  std_logic_vector(46 downto 0);
   -- timing of level3: (c10, 0.116154ns)
signal count2, count2_d1 :  std_logic;
   -- timing of count2: (c10, 0.676154ns)
signal level2, level2_d1 :  std_logic_vector(42 downto 0);
   -- timing of level2: (c10, 1.226154ns)
signal count1, count1_d1 :  std_logic;
   -- timing of count1: (c10, 1.786154ns)
signal level1 :  std_logic_vector(40 downto 0);
   -- timing of level1: (c11, 0.536154ns)
signal count0 :  std_logic;
   -- timing of count0: (c11, 1.096154ns)
signal level0 :  std_logic_vector(39 downto 0);
   -- timing of level0: (c11, 1.646154ns)
signal sCount :  std_logic_vector(4 downto 0);
   -- timing of sCount: (c11, 1.096154ns)
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            level5_d1 <=  level5;
            count4_d1 <=  count4;
            count4_d2 <=  count4_d1;
            level4_d1 <=  level4;
            count3_d1 <=  count3;
            count3_d2 <=  count3_d1;
            count2_d1 <=  count2;
            level2_d1 <=  level2;
            count1_d1 <=  count1;
         end if;
      end process;
   level5 <= X ;
   count4<= '1' when level5_d1(47 downto 32) = (47 downto 32=>'0') else '0';
   level4<= level5_d1(47 downto 0) when count4='0' else level5_d1(31 downto 0) & (15 downto 0 => '0');

   count3<= '1' when level4(47 downto 40) = (47 downto 40=>'0') else '0';
   level3<= level4_d1(47 downto 1) when count3_d1='0' else level4_d1(39 downto 0) & (6 downto 0 => '0');

   count2<= '1' when level3(46 downto 43) = (46 downto 43=>'0') else '0';
   level2<= level3(46 downto 4) when count2='0' else level3(42 downto 0);

   count1<= '1' when level2(42 downto 41) = (42 downto 41=>'0') else '0';
   level1<= level2_d1(42 downto 2) when count1_d1='0' else level2_d1(40 downto 0);

   count0<= '1' when level1(40 downto 40) = (40 downto 40=>'0') else '0';
   level0<= level1(40 downto 1) when count0='0' else level1(39 downto 0);

   R <= level0;
   sCount <= count4_d2 & count3_d2 & count2_d1 & count1_d1 & count0;
   Count <= sCount;
end architecture;

--------------------------------------------------------------------------------
--                   RightShifter16_by_max_15_Freq500_uid47
-- VHDL generated for DummyFPGA @ 500MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca (2008-2011), Florent de Dinechin (2008-2019)
--------------------------------------------------------------------------------
-- Pipeline depth: 3 cycles
-- Clock period (ns): 2
-- Target frequency (MHz): 500
-- Input signals: X S
-- Output signals: R
--  approx. input signal timings: X: (c5, 0.156154ns)S: (c3, 1.460000ns)
--  approx. output signal timings: R: (c6, 0.225385ns)

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity RightShifter16_by_max_15_Freq500_uid47 is
    port (clk : in std_logic;
          X : in  std_logic_vector(15 downto 0);
          S : in  std_logic_vector(3 downto 0);
          R : out  std_logic_vector(30 downto 0)   );
end entity;

architecture arch of RightShifter16_by_max_15_Freq500_uid47 is
signal ps, ps_d1, ps_d2, ps_d3 :  std_logic_vector(3 downto 0);
   -- timing of ps: (c3, 1.460000ns)
signal level0 :  std_logic_vector(15 downto 0);
   -- timing of level0: (c5, 0.156154ns)
signal level1 :  std_logic_vector(16 downto 0);
   -- timing of level1: (c5, 0.156154ns)
signal level2 :  std_logic_vector(18 downto 0);
   -- timing of level2: (c5, 0.998462ns)
signal level3, level3_d1 :  std_logic_vector(22 downto 0);
   -- timing of level3: (c5, 0.998462ns)
signal level4 :  std_logic_vector(30 downto 0);
   -- timing of level4: (c6, 0.225385ns)
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            ps_d1 <=  ps;
            ps_d2 <=  ps_d1;
            ps_d3 <=  ps_d2;
            level3_d1 <=  level3;
         end if;
      end process;
   ps<= S;
   level0<= X;
   level1 <=  (0 downto 0 => '0') & level0 when ps_d2(0) = '1' else    level0 & (0 downto 0 => '0');
   level2 <=  (1 downto 0 => '0') & level1 when ps_d2(1) = '1' else    level1 & (1 downto 0 => '0');
   level3 <=  (3 downto 0 => '0') & level2 when ps_d2(2) = '1' else    level2 & (3 downto 0 => '0');
   level4 <=  (7 downto 0 => '0') & level3_d1 when ps_d3(3) = '1' else    level3_d1 & (7 downto 0 => '0');
   R <= level4(30 downto 0);
end architecture;

--------------------------------------------------------------------------------
--                         IntAdder_29_Freq500_uid49
-- VHDL generated for DummyFPGA @ 500MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin (2008-2016)
--------------------------------------------------------------------------------
-- Pipeline depth: 6 cycles
-- Clock period (ns): 2
-- Target frequency (MHz): 500
-- Input signals: X Y Cin
-- Output signals: R
--  approx. input signal timings: X: (c4, 1.406154ns)Y: (c6, 0.225385ns)Cin: (c0, 0.550000ns)
--  approx. output signal timings: R: (c6, 1.505385ns)

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntAdder_29_Freq500_uid49 is
    port (clk : in std_logic;
          X : in  std_logic_vector(28 downto 0);
          Y : in  std_logic_vector(28 downto 0);
          Cin : in  std_logic;
          R : out  std_logic_vector(28 downto 0)   );
end entity;

architecture arch of IntAdder_29_Freq500_uid49 is
signal Rtmp :  std_logic_vector(28 downto 0);
   -- timing of Rtmp: (c6, 1.505385ns)
signal X_d1, X_d2 :  std_logic_vector(28 downto 0);
   -- timing of X: (c4, 1.406154ns)
signal Cin_d1, Cin_d2, Cin_d3, Cin_d4, Cin_d5, Cin_d6 :  std_logic;
   -- timing of Cin: (c0, 0.550000ns)
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            X_d1 <=  X;
            X_d2 <=  X_d1;
            Cin_d1 <=  Cin;
            Cin_d2 <=  Cin_d1;
            Cin_d3 <=  Cin_d2;
            Cin_d4 <=  Cin_d3;
            Cin_d5 <=  Cin_d4;
            Cin_d6 <=  Cin_d5;
         end if;
      end process;
   Rtmp <= X_d2 + Y + Cin_d6;
   R <= Rtmp;
end architecture;

--------------------------------------------------------------------------------
--                         IntAdder_31_Freq500_uid52
-- VHDL generated for DummyFPGA @ 500MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin (2008-2016)
--------------------------------------------------------------------------------
-- Pipeline depth: 12 cycles
-- Clock period (ns): 2
-- Target frequency (MHz): 500
-- Input signals: X Y Cin
-- Output signals: R
--  approx. input signal timings: X: (c11, 1.646154ns)Y: (c11, 1.646154ns)Cin: (c0, 0.000000ns)
--  approx. output signal timings: R: (c12, 1.156154ns)

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntAdder_31_Freq500_uid52 is
    port (clk : in std_logic;
          X : in  std_logic_vector(30 downto 0);
          Y : in  std_logic_vector(30 downto 0);
          Cin : in  std_logic;
          R : out  std_logic_vector(30 downto 0)   );
end entity;

architecture arch of IntAdder_31_Freq500_uid52 is
signal Cin_1, Cin_1_d1, Cin_1_d2, Cin_1_d3, Cin_1_d4, Cin_1_d5, Cin_1_d6, Cin_1_d7, Cin_1_d8, Cin_1_d9, Cin_1_d10, Cin_1_d11, Cin_1_d12 :  std_logic;
   -- timing of Cin_1: (c0, 0.000000ns)
signal X_1, X_1_d1 :  std_logic_vector(31 downto 0);
   -- timing of X_1: (c11, 1.646154ns)
signal Y_1, Y_1_d1 :  std_logic_vector(31 downto 0);
   -- timing of Y_1: (c11, 1.646154ns)
signal S_1 :  std_logic_vector(31 downto 0);
   -- timing of S_1: (c12, 1.156154ns)
signal R_1 :  std_logic_vector(30 downto 0);
   -- timing of R_1: (c12, 1.156154ns)
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            Cin_1_d1 <=  Cin_1;
            Cin_1_d2 <=  Cin_1_d1;
            Cin_1_d3 <=  Cin_1_d2;
            Cin_1_d4 <=  Cin_1_d3;
            Cin_1_d5 <=  Cin_1_d4;
            Cin_1_d6 <=  Cin_1_d5;
            Cin_1_d7 <=  Cin_1_d6;
            Cin_1_d8 <=  Cin_1_d7;
            Cin_1_d9 <=  Cin_1_d8;
            Cin_1_d10 <=  Cin_1_d9;
            Cin_1_d11 <=  Cin_1_d10;
            Cin_1_d12 <=  Cin_1_d11;
            X_1_d1 <=  X_1;
            Y_1_d1 <=  Y_1;
         end if;
      end process;
   Cin_1 <= Cin;
   X_1 <= '0' & X(30 downto 0);
   Y_1 <= '0' & Y(30 downto 0);
   S_1 <= X_1_d1 + Y_1_d1 + Cin_1_d12;
   R_1 <= S_1(30 downto 0);
   R <= R_1 ;
end architecture;

--------------------------------------------------------------------------------
--                                 top_module
--                  (FPLogIterative_8_23_0_500_Freq500_uid2)
-- VHDL generated for DummyFPGA @ 500MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: F. de Dinechin, C. Klein  (2008-2011)
--------------------------------------------------------------------------------
-- Pipeline depth: 12 cycles
-- Clock period (ns): 2
-- Target frequency (MHz): 500
-- Input signals: X
-- Output signals: R
--  approx. input signal timings: X: (c0, 0.000000ns)
--  approx. output signal timings: R: (c12, 1.156154ns)

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity top_module is
    port (clk : in std_logic;
          X : in  std_logic_vector(8+23+2 downto 0);
          R : out  std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of top_module is
   component LZOC_23_Freq500_uid4 is
      port ( clk : in std_logic;
             I : in  std_logic_vector(22 downto 0);
             OZB : in  std_logic;
             O : out  std_logic_vector(4 downto 0)   );
   end component;

   component LeftShifter12_by_max_12_Freq500_uid6 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(11 downto 0);
             S : in  std_logic_vector(3 downto 0);
             R : out  std_logic_vector(23 downto 0)   );
   end component;

   component InvA0Table_Freq500_uid8 is
      port ( X : in  std_logic_vector(8 downto 0);
             Y : out  std_logic_vector(9 downto 0)   );
   end component;

   component IntAdder_27_Freq500_uid12 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(26 downto 0);
             Y : in  std_logic_vector(26 downto 0);
             Cin : in  std_logic;
             R : out  std_logic_vector(26 downto 0)   );
   end component;

   component IntAdder_27_Freq500_uid15 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(26 downto 0);
             Y : in  std_logic_vector(26 downto 0);
             Cin : in  std_logic;
             R : out  std_logic_vector(26 downto 0)   );
   end component;

   component IntAdder_27_Freq500_uid18 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(26 downto 0);
             Y : in  std_logic_vector(26 downto 0);
             Cin : in  std_logic;
             R : out  std_logic_vector(26 downto 0)   );
   end component;

   component LogTable0_Freq500_uid20 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(8 downto 0);
             Y : out  std_logic_vector(39 downto 0)   );
   end component;

   component LogTable1_Freq500_uid22 is
      port ( X : in  std_logic_vector(6 downto 0);
             Y : out  std_logic_vector(32 downto 0)   );
   end component;

   component IntAdder_40_Freq500_uid26 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(39 downto 0);
             Y : in  std_logic_vector(39 downto 0);
             Cin : in  std_logic;
             R : out  std_logic_vector(39 downto 0)   );
   end component;

   component IntAdder_40_Freq500_uid29 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(39 downto 0);
             Y : in  std_logic_vector(39 downto 0);
             Cin : in  std_logic;
             R : out  std_logic_vector(39 downto 0)   );
   end component;

   component FixRealKCM_Freq500_uid31 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(7 downto 0);
             R : out  std_logic_vector(34 downto 0)   );
   end component;

   component IntAdder_48_Freq500_uid43 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(47 downto 0);
             Y : in  std_logic_vector(47 downto 0);
             Cin : in  std_logic;
             R : out  std_logic_vector(47 downto 0)   );
   end component;

   component Normalizer_Z_48_40_19_Freq500_uid45 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(47 downto 0);
             Count : out  std_logic_vector(4 downto 0);
             R : out  std_logic_vector(39 downto 0)   );
   end component;

   component RightShifter16_by_max_15_Freq500_uid47 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(15 downto 0);
             S : in  std_logic_vector(3 downto 0);
             R : out  std_logic_vector(30 downto 0)   );
   end component;

   component IntAdder_29_Freq500_uid49 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(28 downto 0);
             Y : in  std_logic_vector(28 downto 0);
             Cin : in  std_logic;
             R : out  std_logic_vector(28 downto 0)   );
   end component;

   component IntAdder_31_Freq500_uid52 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(30 downto 0);
             Y : in  std_logic_vector(30 downto 0);
             Cin : in  std_logic;
             R : out  std_logic_vector(30 downto 0)   );
   end component;

signal XExnSgn, XExnSgn_d1, XExnSgn_d2, XExnSgn_d3, XExnSgn_d4, XExnSgn_d5, XExnSgn_d6, XExnSgn_d7, XExnSgn_d8, XExnSgn_d9, XExnSgn_d10, XExnSgn_d11, XExnSgn_d12 :  std_logic_vector(2 downto 0);
   -- timing of XExnSgn: (c0, 0.000000ns)
signal FirstBit :  std_logic;
   -- timing of FirstBit: (c0, 0.000000ns)
signal Y0, Y0_d1 :  std_logic_vector(24 downto 0);
   -- timing of Y0: (c0, 0.550000ns)
signal Y0h :  std_logic_vector(22 downto 0);
   -- timing of Y0h: (c0, 0.550000ns)
signal sR, sR_d1, sR_d2, sR_d3, sR_d4, sR_d5, sR_d6, sR_d7, sR_d8, sR_d9, sR_d10, sR_d11, sR_d12 :  std_logic;
   -- timing of sR: (c0, 0.550000ns)
signal absZ0 :  std_logic_vector(11 downto 0);
   -- timing of absZ0: (c0, 1.660000ns)
signal E :  std_logic_vector(7 downto 0);
   -- timing of E: (c0, 1.070000ns)
signal absE :  std_logic_vector(7 downto 0);
   -- timing of absE: (c0, 1.620000ns)
signal EeqZero, EeqZero_d1, EeqZero_d2, EeqZero_d3, EeqZero_d4 :  std_logic;
   -- timing of EeqZero: (c0, 1.620000ns)
signal lzo, lzo_d1, lzo_d2, lzo_d3 :  std_logic_vector(4 downto 0);
   -- timing of lzo: (c3, 0.410000ns)
signal pfinal_s, pfinal_s_d1, pfinal_s_d2, pfinal_s_d3 :  std_logic_vector(4 downto 0);
   -- timing of pfinal_s: (c0, 0.000000ns)
signal shiftval :  std_logic_vector(5 downto 0);
   -- timing of shiftval: (c3, 1.460000ns)
signal shiftvalinL :  std_logic_vector(3 downto 0);
   -- timing of shiftvalinL: (c3, 1.460000ns)
signal shiftvalinR :  std_logic_vector(3 downto 0);
   -- timing of shiftvalinR: (c3, 1.460000ns)
signal doRR, doRR_d1, doRR_d2 :  std_logic;
   -- timing of doRR: (c3, 1.460000ns)
signal small, small_d1, small_d2, small_d3, small_d4, small_d5, small_d6, small_d7, small_d8 :  std_logic;
   -- timing of small: (c4, 0.210000ns)
signal small_absZ0_normd_full :  std_logic_vector(23 downto 0);
   -- timing of small_absZ0_normd_full: (c4, 1.406154ns)
signal small_absZ0_normd, small_absZ0_normd_d1 :  std_logic_vector(11 downto 0);
   -- timing of small_absZ0_normd: (c4, 1.406154ns)
signal A0 :  std_logic_vector(8 downto 0);
   -- timing of A0: (c0, 0.000000ns)
signal InvA0, InvA0_d1 :  std_logic_vector(9 downto 0);
   -- timing of InvA0: (c0, 0.550000ns)
signal InvA0_copy9 :  std_logic_vector(9 downto 0);
   -- timing of InvA0_copy9: (c0, 0.000000ns)
signal P0 :  std_logic_vector(34 downto 0);
   -- timing of P0: (c1, 0.640000ns)
signal Z1 :  std_logic_vector(25 downto 0);
   -- timing of Z1: (c1, 0.640000ns)
signal A1, A1_d1 :  std_logic_vector(6 downto 0);
   -- timing of A1: (c1, 0.640000ns)
signal B1 :  std_logic_vector(18 downto 0);
   -- timing of B1: (c1, 0.640000ns)
signal ZM1, ZM1_d1 :  std_logic_vector(25 downto 0);
   -- timing of ZM1: (c1, 0.640000ns)
signal P1 :  std_logic_vector(32 downto 0);
   -- timing of P1: (c2, 0.710000ns)
signal Y1 :  std_logic_vector(33 downto 0);
   -- timing of Y1: (c1, 0.640000ns)
signal EiY1 :  std_logic_vector(26 downto 0);
   -- timing of EiY1: (c1, 1.190000ns)
signal addXIter1 :  std_logic_vector(26 downto 0);
   -- timing of addXIter1: (c1, 0.640000ns)
signal EiYPB1 :  std_logic_vector(26 downto 0);
   -- timing of EiYPB1: (c2, 0.660000ns)
signal Pp1 :  std_logic_vector(26 downto 0);
   -- timing of Pp1: (c2, 1.260000ns)
signal Z2 :  std_logic_vector(26 downto 0);
   -- timing of Z2: (c3, 0.730000ns)
signal Zfinal, Zfinal_d1, Zfinal_d2 :  std_logic_vector(26 downto 0);
   -- timing of Zfinal: (c3, 0.730000ns)
signal squarerIn :  std_logic_vector(15 downto 0);
   -- timing of squarerIn: (c5, 0.156154ns)
signal Z2o2_full :  std_logic_vector(31 downto 0);
   -- timing of Z2o2_full: (c5, 0.156154ns)
signal Z2o2_full_dummy :  std_logic_vector(31 downto 0);
   -- timing of Z2o2_full_dummy: (c5, 0.156154ns)
signal Z2o2_normal :  std_logic_vector(12 downto 0);
   -- timing of Z2o2_normal: (c5, 0.156154ns)
signal addFinalLog1pY :  std_logic_vector(26 downto 0);
   -- timing of addFinalLog1pY: (c5, 0.706154ns)
signal Log1p_normal :  std_logic_vector(26 downto 0);
   -- timing of Log1p_normal: (c6, 1.176154ns)
signal L0 :  std_logic_vector(39 downto 0);
   -- timing of L0: (c2, 0.415625ns)
signal S1 :  std_logic_vector(39 downto 0);
   -- timing of S1: (c2, 0.415625ns)
signal L1 :  std_logic_vector(32 downto 0);
   -- timing of L1: (c1, 1.190000ns)
signal L1_copy23 :  std_logic_vector(32 downto 0);
   -- timing of L1_copy23: (c1, 0.640000ns)
signal sopX1 :  std_logic_vector(39 downto 0);
   -- timing of sopX1: (c1, 1.190000ns)
signal S2 :  std_logic_vector(39 downto 0);
   -- timing of S2: (c3, 1.015625ns)
signal almostLog :  std_logic_vector(39 downto 0);
   -- timing of almostLog: (c3, 1.015625ns)
signal adderLogF_normalY :  std_logic_vector(39 downto 0);
   -- timing of adderLogF_normalY: (c6, 1.176154ns)
signal LogF_normal :  std_logic_vector(39 downto 0);
   -- timing of LogF_normal: (c7, 0.776154ns)
signal absELog2 :  std_logic_vector(34 downto 0);
   -- timing of absELog2: (c1, 1.710000ns)
signal absELog2_pad :  std_logic_vector(47 downto 0);
   -- timing of absELog2_pad: (c1, 1.710000ns)
signal LogF_normal_pad :  std_logic_vector(47 downto 0);
   -- timing of LogF_normal_pad: (c7, 0.776154ns)
signal lnaddX :  std_logic_vector(47 downto 0);
   -- timing of lnaddX: (c1, 1.710000ns)
signal lnaddY :  std_logic_vector(47 downto 0);
   -- timing of lnaddY: (c7, 0.776154ns)
signal Log_normal :  std_logic_vector(47 downto 0);
   -- timing of Log_normal: (c8, 1.456154ns)
signal Log_normal_normd, Log_normal_normd_d1 :  std_logic_vector(39 downto 0);
   -- timing of Log_normal_normd: (c11, 1.646154ns)
signal E_normal :  std_logic_vector(4 downto 0);
   -- timing of E_normal: (c11, 1.096154ns)
signal Z2o2_small_bs :  std_logic_vector(15 downto 0);
   -- timing of Z2o2_small_bs: (c5, 0.156154ns)
signal Z2o2_small_s :  std_logic_vector(30 downto 0);
   -- timing of Z2o2_small_s: (c6, 0.225385ns)
signal Z2o2_small :  std_logic_vector(28 downto 0);
   -- timing of Z2o2_small: (c6, 0.225385ns)
signal Z_small :  std_logic_vector(28 downto 0);
   -- timing of Z_small: (c4, 1.406154ns)
signal Log_smallY :  std_logic_vector(28 downto 0);
   -- timing of Log_smallY: (c6, 0.225385ns)
signal nsRCin :  std_logic;
   -- timing of nsRCin: (c0, 0.550000ns)
signal Log_small :  std_logic_vector(28 downto 0);
   -- timing of Log_small: (c6, 1.505385ns)
signal E0_sub :  std_logic_vector(1 downto 0);
   -- timing of E0_sub: (c6, 1.505385ns)
signal ufl, ufl_d1, ufl_d2, ufl_d3, ufl_d4, ufl_d5, ufl_d6, ufl_d7, ufl_d8, ufl_d9, ufl_d10, ufl_d11, ufl_d12 :  std_logic;
   -- timing of ufl: (c0, 0.000000ns)
signal E_small, E_small_d1, E_small_d2, E_small_d3, E_small_d4, E_small_d5 :  std_logic_vector(7 downto 0);
   -- timing of E_small: (c6, 1.505385ns)
signal Log_small_normd, Log_small_normd_d1, Log_small_normd_d2, Log_small_normd_d3, Log_small_normd_d4, Log_small_normd_d5, Log_small_normd_d6 :  std_logic_vector(26 downto 0);
   -- timing of Log_small_normd: (c6, 1.505385ns)
signal E0offset, E0offset_d1, E0offset_d2, E0offset_d3, E0offset_d4, E0offset_d5, E0offset_d6, E0offset_d7, E0offset_d8, E0offset_d9, E0offset_d10, E0offset_d11 :  std_logic_vector(7 downto 0);
   -- timing of E0offset: (c0, 0.000000ns)
signal ER :  std_logic_vector(7 downto 0);
   -- timing of ER: (c11, 1.096154ns)
signal Log_g :  std_logic_vector(26 downto 0);
   -- timing of Log_g: (c11, 1.646154ns)
signal round :  std_logic;
   -- timing of round: (c11, 1.646154ns)
signal fraX :  std_logic_vector(30 downto 0);
   -- timing of fraX: (c11, 1.646154ns)
signal fraY :  std_logic_vector(30 downto 0);
   -- timing of fraY: (c11, 1.646154ns)
signal EFR :  std_logic_vector(30 downto 0);
   -- timing of EFR: (c12, 1.156154ns)
signal Rexn :  std_logic_vector(2 downto 0);
   -- timing of Rexn: (c12, 0.396154ns)
constant g: positive := 4;
constant log2wF: positive := 5;
constant pfinal: positive := 13;
constant sfinal: positive := 27;
constant targetprec: positive := 40;
constant wE: positive := 8;
constant wF: positive := 23;
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            XExnSgn_d1 <=  XExnSgn;
            XExnSgn_d2 <=  XExnSgn_d1;
            XExnSgn_d3 <=  XExnSgn_d2;
            XExnSgn_d4 <=  XExnSgn_d3;
            XExnSgn_d5 <=  XExnSgn_d4;
            XExnSgn_d6 <=  XExnSgn_d5;
            XExnSgn_d7 <=  XExnSgn_d6;
            XExnSgn_d8 <=  XExnSgn_d7;
            XExnSgn_d9 <=  XExnSgn_d8;
            XExnSgn_d10 <=  XExnSgn_d9;
            XExnSgn_d11 <=  XExnSgn_d10;
            XExnSgn_d12 <=  XExnSgn_d11;
            Y0_d1 <=  Y0;
            sR_d1 <=  sR;
            sR_d2 <=  sR_d1;
            sR_d3 <=  sR_d2;
            sR_d4 <=  sR_d3;
            sR_d5 <=  sR_d4;
            sR_d6 <=  sR_d5;
            sR_d7 <=  sR_d6;
            sR_d8 <=  sR_d7;
            sR_d9 <=  sR_d8;
            sR_d10 <=  sR_d9;
            sR_d11 <=  sR_d10;
            sR_d12 <=  sR_d11;
            EeqZero_d1 <=  EeqZero;
            EeqZero_d2 <=  EeqZero_d1;
            EeqZero_d3 <=  EeqZero_d2;
            EeqZero_d4 <=  EeqZero_d3;
            lzo_d1 <=  lzo;
            lzo_d2 <=  lzo_d1;
            lzo_d3 <=  lzo_d2;
            pfinal_s_d1 <=  pfinal_s;
            pfinal_s_d2 <=  pfinal_s_d1;
            pfinal_s_d3 <=  pfinal_s_d2;
            doRR_d1 <=  doRR;
            doRR_d2 <=  doRR_d1;
            small_d1 <=  small;
            small_d2 <=  small_d1;
            small_d3 <=  small_d2;
            small_d4 <=  small_d3;
            small_d5 <=  small_d4;
            small_d6 <=  small_d5;
            small_d7 <=  small_d6;
            small_d8 <=  small_d7;
            small_absZ0_normd_d1 <=  small_absZ0_normd;
            InvA0_d1 <=  InvA0;
            A1_d1 <=  A1;
            ZM1_d1 <=  ZM1;
            Zfinal_d1 <=  Zfinal;
            Zfinal_d2 <=  Zfinal_d1;
            Log_normal_normd_d1 <=  Log_normal_normd;
            ufl_d1 <=  ufl;
            ufl_d2 <=  ufl_d1;
            ufl_d3 <=  ufl_d2;
            ufl_d4 <=  ufl_d3;
            ufl_d5 <=  ufl_d4;
            ufl_d6 <=  ufl_d5;
            ufl_d7 <=  ufl_d6;
            ufl_d8 <=  ufl_d7;
            ufl_d9 <=  ufl_d8;
            ufl_d10 <=  ufl_d9;
            ufl_d11 <=  ufl_d10;
            ufl_d12 <=  ufl_d11;
            E_small_d1 <=  E_small;
            E_small_d2 <=  E_small_d1;
            E_small_d3 <=  E_small_d2;
            E_small_d4 <=  E_small_d3;
            E_small_d5 <=  E_small_d4;
            Log_small_normd_d1 <=  Log_small_normd;
            Log_small_normd_d2 <=  Log_small_normd_d1;
            Log_small_normd_d3 <=  Log_small_normd_d2;
            Log_small_normd_d4 <=  Log_small_normd_d3;
            Log_small_normd_d5 <=  Log_small_normd_d4;
            Log_small_normd_d6 <=  Log_small_normd_d5;
            E0offset_d1 <=  E0offset;
            E0offset_d2 <=  E0offset_d1;
            E0offset_d3 <=  E0offset_d2;
            E0offset_d4 <=  E0offset_d3;
            E0offset_d5 <=  E0offset_d4;
            E0offset_d6 <=  E0offset_d5;
            E0offset_d7 <=  E0offset_d6;
            E0offset_d8 <=  E0offset_d7;
            E0offset_d9 <=  E0offset_d8;
            E0offset_d10 <=  E0offset_d9;
            E0offset_d11 <=  E0offset_d10;
         end if;
      end process;
   XExnSgn <=  X(wE+wF+2 downto wE+wF);
   FirstBit <=  X(wF-1);
   Y0 <= "1" & X(wF-1 downto 0) & "0" when FirstBit = '0' else "01" & X(wF-1 downto 0);
   Y0h <= Y0(wF downto 1);
   -- Sign of the result;
   sR <= '0'   when  (X(wE+wF-1 downto wF) = ('0' & (wE-2 downto 0 => '1')))  -- binade [1..2)
     else not X(wE+wF-1);                -- MSB of exponent
   absZ0 <=   Y0(wF-pfinal+1 downto 0)          when (sR='0') else
             ((wF-pfinal+1 downto 0 => '0') - Y0(wF-pfinal+1 downto 0));
   E <= (X(wE+wF-1 downto wF)) - ("0" & (wE-2 downto 1 => '1') & (not FirstBit));
   absE <= ((wE-1 downto 0 => '0') - E)   when sR = '1' else E;
   EeqZero <= '1' when E=(wE-1 downto 0 => '0') else '0';
   lzoc1: LZOC_23_Freq500_uid4
      port map ( clk  => clk,
                 I => Y0h,
                 OZB => FirstBit,
                 O => lzo);
   pfinal_s <= "01101";
   shiftval <= ('0' & lzo) - ('0' & pfinal_s_d3); 
   shiftvalinL <= shiftval(3 downto 0);
   shiftvalinR <= shiftval(3 downto 0);
   doRR <= shiftval(log2wF); -- sign of the result
   small <= EeqZero_d4 and not(doRR_d1);
   -- The left shifter for the 'small' case
   small_lshift: LeftShifter12_by_max_12_Freq500_uid6
      port map ( clk  => clk,
                 S => shiftvalinL,
                 X => absZ0,
                 R => small_absZ0_normd_full);
   small_absZ0_normd <= small_absZ0_normd_full(11 downto 0); -- get rid of leading zeroes
   ---------------- The range reduction box ---------------
   A0 <= X(22 downto 14);
   -- First inv table
   InvA0Table: InvA0Table_Freq500_uid8
      port map ( X => A0,
                 Y => InvA0_copy9);
   InvA0 <= InvA0_copy9; -- output copy to hold a pipeline register if needed
   P0 <= InvA0_d1 * Y0_d1;

   Z1 <= P0(25 downto 0);

   A1 <= Z1(25 downto 19);
   B1 <= Z1(18 downto 0);
   ZM1 <= Z1;
   P1 <= A1_d1*ZM1_d1;
   Y1 <= "1" & (6 downto 0 => '0') & Z1;
   EiY1 <= Y1(33 downto 7)  when A1(6) = '1'
     else  "0" & Y1(33 downto 8);
   addXIter1 <= "0" & B1 & (6 downto 0 => '0');
   addIter1_1: IntAdder_27_Freq500_uid12
      port map ( clk  => clk,
                 Cin => '0',
                 X => addXIter1,
                 Y => EiY1,
                 R => EiYPB1);
   Pp1 <= (0 downto 0 => '1') & not(P1(32 downto 7));
   addIter2_1: IntAdder_27_Freq500_uid15
      port map ( clk  => clk,
                 Cin => '1',
                 X => EiYPB1,
                 Y => Pp1,
                 R => Z2);
   Zfinal <= Z2;
   squarerIn <= Zfinal_d2(sfinal-1 downto sfinal-16) when doRR_d2='1'
                    else (small_absZ0_normd_d1 & (3 downto 0 => '0'));  
   Z2o2_full <= squarerIn*squarerIn;
   Z2o2_full_dummy <= Z2o2_full;
   Z2o2_normal <= Z2o2_full_dummy (31  downto 19);
   addFinalLog1pY <= (pfinal downto 0  => '1') & not(Z2o2_normal);
   addFinalLog1p_normalAdder: IntAdder_27_Freq500_uid18
      port map ( clk  => clk,
                 Cin => '1',
                 X => Zfinal,
                 Y => addFinalLog1pY,
                 R => Log1p_normal);

   -- Now the log tables, as late as possible
   LogTable0: LogTable0_Freq500_uid20
      port map ( clk  => clk,
                 X => A0,
                 Y => L0);
   S1 <= L0;
   LogTable1: LogTable1_Freq500_uid22
      port map ( X => A1,
                 Y => L1_copy23);
   L1 <= L1_copy23; -- output copy to hold a pipeline register if needed
   sopX1 <= ((39 downto 33 => '0') & L1);
   adderS1: IntAdder_40_Freq500_uid26
      port map ( clk  => clk,
                 Cin => '0',
                 X => S1,
                 Y => sopX1,
                 R => S2);
   almostLog <= S2;
   adderLogF_normalY <= ((targetprec-1 downto sfinal => '0') & Log1p_normal);
   adderLogF_normal: IntAdder_40_Freq500_uid29
      port map ( clk  => clk,
                 Cin => '0',
                 X => almostLog,
                 Y => adderLogF_normalY,
                 R => LogF_normal);
   MulLog2: FixRealKCM_Freq500_uid31
      port map ( clk  => clk,
                 X => absE,
                 R => absELog2);
   absELog2_pad <=   absELog2 & (targetprec-wF-g-1 downto 0 => '0');       
   LogF_normal_pad <= (wE-1  downto 0 => LogF_normal(targetprec-1))  & LogF_normal;
   lnaddX <= absELog2_pad;
   lnaddY <= LogF_normal_pad when sR_d7='0' else not(LogF_normal_pad); 
   lnadder: IntAdder_48_Freq500_uid43
      port map ( clk  => clk,
                 Cin => sR,
                 X => lnaddX,
                 Y => lnaddY,
                 R => Log_normal);
   final_norm: Normalizer_Z_48_40_19_Freq500_uid45
      port map ( clk  => clk,
                 X => Log_normal,
                 Count => E_normal,
                 R => Log_normal_normd);
   Z2o2_small_bs <= Z2o2_full_dummy(31 downto 16);
   ao_rshift: RightShifter16_by_max_15_Freq500_uid47
      port map ( clk  => clk,
                 S => shiftvalinR,
                 X => Z2o2_small_bs,
                 R => Z2o2_small_s);
     -- send the MSB to position pfinal
   Z2o2_small <=  (pfinal-1 downto 0  => '0') & Z2o2_small_s(30 downto 15);
   -- mantissa will be either Y0-z^2/2  or  -Y0+z^2/2,  depending on sR  
   Z_small <= small_absZ0_normd & (16 downto 0 => '0');
   Log_smallY <= Z2o2_small when sR_d6='1' else not(Z2o2_small);
   nsRCin <= not ( sR );
   log_small_adder: IntAdder_29_Freq500_uid49
      port map ( clk  => clk,
                 Cin => nsRCin,
                 X => Z_small,
                 Y => Log_smallY,
                 R => Log_small);
   -- Possibly subtract 1 or 2 to the exponent, depending on the LZC of Log_small
   E0_sub <=   "11" when Log_small(wF+g+1) = '1'
          else "10" when Log_small(wF+g+1 downto wF+g) = "01"
          else "01" ;
   -- The smallest log will be log(1+2^{-wF}) \approx 2^{-wF}  = 2^-23
   -- The smallest representable number is 2^{1-2^(wE-1)} = 2^-127
   -- No underflow possible
   ufl <= '0';
   E_small <=  ("0" & (wE-2 downto 2 => '1') & E0_sub)  -  ((wE-1 downto 5 => '0') & lzo_d3) ;
   Log_small_normd <= Log_small(wF+g+1 downto 2) when Log_small(wF+g+1)='1'
           else Log_small(wF+g downto 1)  when Log_small(wF+g)='1'  -- remove the first zero
           else Log_small(wF+g-1 downto 0)  ; -- remove two zeroes (extremely rare, 001000000 only)
   E0offset <= "10000110"; -- E0 + wE 
   ER <= E_small_d5(7 downto 0) when small_d7='1'
      else E0offset_d11 - ((7 downto 5 => '0') & E_normal);
   Log_g <=  Log_small_normd_d5(wF+g-2 downto 0) & "0" when small_d7='1'           -- remove implicit 1
      else Log_normal_normd(targetprec-2 downto targetprec-wF-g-1 );  -- remove implicit 1
   round <= Log_g(g-1) ; -- sticky is always 1 for a transcendental function 
   -- if round leads to a change of binade, the carry propagation magically updates both mantissa and exponent
   fraX <= (ER & Log_g(wF+g-1 downto g)) ; 
   fraY <= ((wE+wF-1 downto 1 => '0') & round); 
   finalRoundAdder: IntAdder_31_Freq500_uid52
      port map ( clk  => clk,
                 Cin => '0',
                 X => fraX,
                 Y => fraY,
                 R => EFR);
   Rexn <= "110" when ((XExnSgn_d12(2) and (XExnSgn_d12(1) or XExnSgn_d12(0))) or (XExnSgn_d12(1) and XExnSgn_d12(0))) = '1' else
                              "101" when XExnSgn_d12(2 downto 1) = "00"  else
                              "100" when XExnSgn_d12(2 downto 1) = "10"  else
                              "00" & sR_d12 when (((Log_normal_normd_d1(targetprec-1)='0') and (small_d8='0')) or ( (Log_small_normd_d6 (wF+g-1)='0') and (small_d8='1'))) or (ufl_d12 = '1' and small_d8='1') else
                               "01" & sR_d12;
   R<=  Rexn & EFR;
end architecture;

--------------------------------------------------------------------------------
--                     TestBench_top_module_Freq500_uid54
-- VHDL generated for DummyFPGA @ 500MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Cristian Klein, Nicolas Brunie (2007-2010)
--------------------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity TestBench_top_module_Freq500_uid54 is
end entity;

architecture behavorial of TestBench_top_module_Freq500_uid54 is
   component top_module is
      port ( clk : in std_logic;
             X : in  std_logic_vector(8+23+2 downto 0);
             R : out  std_logic_vector(8+23+2 downto 0)   );
   end component;
signal X :  std_logic_vector(33 downto 0);
   -- timing of X: (c0, 0.000000ns)
signal R :  std_logic_vector(33 downto 0);
   -- timing of R: (c12, 0.000000ns)
signal clk :  std_logic;
   -- timing of clk: (c0, 0.000000ns)
signal rst :  std_logic;
   -- timing of rst: (c0, 0.000000ns)

 -- converts std_logic into a character
   function chr(sl: std_logic) return character is
      variable c: character;
   begin
      case sl is
         when 'U' => c:= 'U';
         when 'X' => c:= 'X';
         when '0' => c:= '0';
         when '1' => c:= '1';
         when 'Z' => c:= 'Z';
         when 'W' => c:= 'W';
         when 'L' => c:= 'L';
         when 'H' => c:= 'H';
         when '-' => c:= '-';
      end case;
      return c;
   end chr;

   -- converts bit to std_logic (1 to 1)
   function to_stdlogic(b : bit) return std_logic is
       variable sl : std_logic;
   begin
      case b is 
         when '0' => sl := '0';
         when '1' => sl := '1';
      end case;
      return sl;
   end to_stdlogic;

   -- converts std_logic into a string (1 to 1)
   function str(sl: std_logic) return string is
    variable s: string(1 to 1);
    begin
      s(1) := chr(sl);
      return s;
   end str;

   -- converts std_logic_vector into a string (binary base)
   -- (this also takes care of the fact that the range of
   --  a string is natural while a std_logic_vector may
   --  have an integer range)
   function str(slv: std_logic_vector) return string is
      variable result : string (1 to slv'length);
      variable r : integer;
   begin
      r := 1;
      for i in slv'range loop
         result(r) := chr(slv(i));
         r := r + 1;
      end loop;
      return result;
   end str;

   -- FP compare function (found vs. real)
   function fp_equal(a : std_logic_vector; b : std_logic_vector) return boolean is
   begin
      if b(b'high downto b'high-1) = "01" then
         return a = b;
      elsif b(b'high downto b'high-1) = "11" then
         return (a(a'high downto a'high-1)=b(b'high downto b'high-1));
      else
         return a(a'high downto a'high-2) = b(b'high downto b'high-2);
      end if;
   end;

   function fp_inf_or_equal(a : std_logic_vector; b : std_logic_vector) return boolean is
   begin
      if (b(b'high downto b'high-1) = "11") or (a(a'high downto a'high-1) = "11")  then
         return false; -- NaN always compare false
      else return true; -- TODO
      end if;
   end;

   -- FP subtypes for casting
   subtype fp34 is std_logic_vector(33 downto 0);
   function testLine(testCounter:integer; expectedOutputS: string(1 to 10000); expectedOutputSize: integer; R:  std_logic_vector(8+23+2 downto 0)) return boolean is
      variable expectedOutput: line;
      variable possibilityNumber : integer;
      variable testSuccess: boolean;
      variable errorMessage: string(1 to 10000);
      variable testSuccess_R: boolean;
      variable expected_R: bit_vector (33 downto 0); -- for list of values
      variable inf_R: bit_vector (33 downto 0); -- for intervals
      variable sup_R: bit_vector (33 downto 0); -- for intervals
   begin
      write(expectedOutput, expectedOutputS);
      read(expectedOutput, possibilityNumber); -- for R
      if possibilityNumber = 0 then
         -- TODO define what it means to have 0 possible output. Currently it means a test fails...
      end if;
      if possibilityNumber > 0 then -- a list of values
      testSuccess_R := false;
         for i in 1 to possibilityNumber loop
            read(expectedOutput, expected_R);
            if fp_equal(R, to_stdlogicvector(expected_R)) then
               testSuccess_R := true;
            end if;
            end loop;
      end if;
      if possibilityNumber < 0  then -- an interval
         read(expectedOutput, inf_R);
         read(expectedOutput, sup_R);
         if possibilityNumber =-1  then -- an unsigned interval
            testSuccess_R := (R >= to_stdlogicvector(inf_R)) and (R <= to_stdlogicvector(sup_R));
         elsif possibilityNumber =-2  then -- a signed interval
            testSuccess_R := (signed(R) >= signed(to_stdlogicvector(inf_R))) and (signed(R) <= signed(to_stdlogicvector(sup_R)));
         elsif possibilityNumber =-4  then -- a floating-point interval
            testSuccess_R := fp_inf_or_equal(to_stdlogicvector(inf_R), R) and fp_inf_or_equal(R, to_stdlogicvector(sup_R));
         end if;
      end if;
      if testSuccess_R = false then
         report("Test #" & integer'image(testCounter) & ", incorrect output for R: " & lf & " expected values: " & expectedOutputS(1 to expectedOutputSize) & lf  & "          result:    " & str(R) ) severity error;
      end if;
      
      testSuccess := true and testSuccess_R;
      return testSuccess;
   end testLine;

begin
   -- Ticking clock signal
   process
   begin
      clk <= '0';
      wait for 5 ns;
      clk <= '1';
      wait for 5 ns;
   end process;

   test: top_module
      port map ( clk  => clk,
                 X => X,
                 R => R);
   -- Process that sets the inputs  (read from a file) 
   process
      variable input, expectedOutput : line; 
      variable tmpChar : character;
      file inputsFile : text is "test.input"; 
      variable V_X : bit_vector(33 downto 0);
      variable V_R : bit_vector(33 downto 0);
   begin
      -- Send reset
      rst <= '1';
      wait for 10 ns;
      rst <= '0';
      readline(inputsFile, input); -- skip the first line of advertising
      while not endfile(inputsFile) loop
         readline(inputsFile, input); -- skip the comment line
         readline(inputsFile, input);
         readline(inputsFile, expectedOutput); -- comment line, unused in this process
         readline(inputsFile, expectedOutput); -- unused in this process
         read(input ,V_X);
         read(input,tmpChar);
         X <= to_stdlogicvector(V_X);
         wait for 10 ns;
      end loop;
         wait for 220 ns; -- wait for pipeline to flush (and some more)
   end process;

    -- Process that verifies the corresponding output
   process
      file inputsFile : text is "test.input"; 
      variable input, expectedOutput : line; 
      variable testCounter : integer := 1;
      variable errorCounter : integer := 0;
      variable expectedOutputString : string(1 to 10000);
      variable testSuccess: boolean;
   begin
      wait for 12 ns; -- wait for reset 
      wait for 120 ns; -- wait for pipeline to flush
      readline(inputsFile, input); -- skip the first line of advertising
      while not endfile(inputsFile) loop
         readline(inputsFile, input); -- input comment, unused
         readline(inputsFile, input); -- input line, unused
         readline(inputsFile, expectedOutput); -- comment line, unused in this process
         readline(inputsFile, expectedOutput);
         expectedOutputString := expectedOutput.all & (expectedOutput'Length+1 to 10000 => ' ');
         testSuccess := testLine(testCounter, expectedOutputString, expectedOutput'Length, R);
         if not testSuccess then 
               errorCounter := errorCounter + 1; -- incrementing global error counter
         end if;
            testCounter := testCounter + 1; -- incrementing global error counter
         wait for 10 ns;
      end loop;
      report integer'image(errorCounter) & " error(s) encoutered." severity note;
      report "End of simulation after " & integer'image(testCounter-1) & " tests" severity note;
   end process;

end architecture;

