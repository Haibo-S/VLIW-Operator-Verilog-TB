module intadder_21_freq500_uid99
  (input  clk,
   input  [20:0] x,
   input  [20:0] y,
   input  cin,
   output [20:0] r);
  wire [20:0] rtmp;
  wire [20:0] x_d1;
  wire [20:0] y_d1;
  wire cin_d1;
  wire cin_d2;
  wire cin_d3;
  wire cin_d4;
  wire cin_d5;
  wire cin_d6;
  wire cin_d7;
  wire cin_d8;
  wire cin_d9;
  wire cin_d10;
  wire cin_d11;
  wire cin_d12;
  wire cin_d13;
  wire cin_d14;
  wire cin_d15;
  wire cin_d16;
  wire cin_d17;
  wire [20:0] n8007;
  wire [20:0] n8008;
  wire [20:0] n8009;
  reg [20:0] n8010;
  reg [20:0] n8011;
  reg n8012;
  reg n8013;
  reg n8014;
  reg n8015;
  reg n8016;
  reg n8017;
  reg n8018;
  reg n8019;
  reg n8020;
  reg n8021;
  reg n8022;
  reg n8023;
  reg n8024;
  reg n8025;
  reg n8026;
  reg n8027;
  reg n8028;
  assign r = rtmp; //(module output)
  /* fppowtf32.vhdl:4669:8  */
  assign rtmp = n8009; // (signal)
  /* fppowtf32.vhdl:4671:8  */
  assign x_d1 = n8010; // (signal)
  /* fppowtf32.vhdl:4673:8  */
  assign y_d1 = n8011; // (signal)
  /* fppowtf32.vhdl:4675:8  */
  assign cin_d1 = n8012; // (signal)
  /* fppowtf32.vhdl:4675:16  */
  assign cin_d2 = n8013; // (signal)
  /* fppowtf32.vhdl:4675:24  */
  assign cin_d3 = n8014; // (signal)
  /* fppowtf32.vhdl:4675:32  */
  assign cin_d4 = n8015; // (signal)
  /* fppowtf32.vhdl:4675:40  */
  assign cin_d5 = n8016; // (signal)
  /* fppowtf32.vhdl:4675:48  */
  assign cin_d6 = n8017; // (signal)
  /* fppowtf32.vhdl:4675:56  */
  assign cin_d7 = n8018; // (signal)
  /* fppowtf32.vhdl:4675:64  */
  assign cin_d8 = n8019; // (signal)
  /* fppowtf32.vhdl:4675:72  */
  assign cin_d9 = n8020; // (signal)
  /* fppowtf32.vhdl:4675:80  */
  assign cin_d10 = n8021; // (signal)
  /* fppowtf32.vhdl:4675:89  */
  assign cin_d11 = n8022; // (signal)
  /* fppowtf32.vhdl:4675:98  */
  assign cin_d12 = n8023; // (signal)
  /* fppowtf32.vhdl:4675:107  */
  assign cin_d13 = n8024; // (signal)
  /* fppowtf32.vhdl:4675:116  */
  assign cin_d14 = n8025; // (signal)
  /* fppowtf32.vhdl:4675:125  */
  assign cin_d15 = n8026; // (signal)
  /* fppowtf32.vhdl:4675:134  */
  assign cin_d16 = n8027; // (signal)
  /* fppowtf32.vhdl:4675:143  */
  assign cin_d17 = n8028; // (signal)
  /* fppowtf32.vhdl:4702:17  */
  assign n8007 = x_d1 + y_d1;
  /* fppowtf32.vhdl:4702:24  */
  assign n8008 = {20'b0, cin_d17};  //  uext
  /* fppowtf32.vhdl:4702:24  */
  assign n8009 = n8007 + n8008;
  /* fppowtf32.vhdl:4680:10  */
  always @(posedge clk)
    n8010 <= x;
  /* fppowtf32.vhdl:4680:10  */
  always @(posedge clk)
    n8011 <= y;
  /* fppowtf32.vhdl:4680:10  */
  always @(posedge clk)
    n8012 <= cin;
  /* fppowtf32.vhdl:4680:10  */
  always @(posedge clk)
    n8013 <= cin_d1;
  /* fppowtf32.vhdl:4680:10  */
  always @(posedge clk)
    n8014 <= cin_d2;
  /* fppowtf32.vhdl:4680:10  */
  always @(posedge clk)
    n8015 <= cin_d3;
  /* fppowtf32.vhdl:4680:10  */
  always @(posedge clk)
    n8016 <= cin_d4;
  /* fppowtf32.vhdl:4680:10  */
  always @(posedge clk)
    n8017 <= cin_d5;
  /* fppowtf32.vhdl:4680:10  */
  always @(posedge clk)
    n8018 <= cin_d6;
  /* fppowtf32.vhdl:4680:10  */
  always @(posedge clk)
    n8019 <= cin_d7;
  /* fppowtf32.vhdl:4680:10  */
  always @(posedge clk)
    n8020 <= cin_d8;
  /* fppowtf32.vhdl:4680:10  */
  always @(posedge clk)
    n8021 <= cin_d9;
  /* fppowtf32.vhdl:4680:10  */
  always @(posedge clk)
    n8022 <= cin_d10;
  /* fppowtf32.vhdl:4680:10  */
  always @(posedge clk)
    n8023 <= cin_d11;
  /* fppowtf32.vhdl:4680:10  */
  always @(posedge clk)
    n8024 <= cin_d12;
  /* fppowtf32.vhdl:4680:10  */
  always @(posedge clk)
    n8025 <= cin_d13;
  /* fppowtf32.vhdl:4680:10  */
  always @(posedge clk)
    n8026 <= cin_d14;
  /* fppowtf32.vhdl:4680:10  */
  always @(posedge clk)
    n8027 <= cin_d15;
  /* fppowtf32.vhdl:4680:10  */
  always @(posedge clk)
    n8028 <= cin_d16;
endmodule

module fixrealkcm_freq500_uid89_t1_freq500_uid95
  (input  [2:0] x,
   output [15:0] y);
  wire [15:0] y0;
  wire [15:0] y1;
  wire n7958;
  wire n7961;
  wire n7964;
  wire n7967;
  wire n7970;
  wire n7973;
  wire n7976;
  wire n7979;
  wire [7:0] n7981;
  reg [15:0] n7982;
  assign y = y1; //(module output)
  /* fppowtf32.vhdl:1062:8  */
  assign y0 = n7982; // (signal)
  /* fppowtf32.vhdl:1064:8  */
  assign y1 = y0; // (signal)
  /* fppowtf32.vhdl:1068:26  */
  assign n7958 = x == 3'b000;
  /* fppowtf32.vhdl:1069:26  */
  assign n7961 = x == 3'b001;
  /* fppowtf32.vhdl:1070:26  */
  assign n7964 = x == 3'b010;
  /* fppowtf32.vhdl:1071:26  */
  assign n7967 = x == 3'b011;
  /* fppowtf32.vhdl:1072:26  */
  assign n7970 = x == 3'b100;
  /* fppowtf32.vhdl:1073:26  */
  assign n7973 = x == 3'b101;
  /* fppowtf32.vhdl:1074:26  */
  assign n7976 = x == 3'b110;
  /* fppowtf32.vhdl:1075:26  */
  assign n7979 = x == 3'b111;
  assign n7981 = {n7979, n7976, n7973, n7970, n7967, n7964, n7961, n7958};
  /* fppowtf32.vhdl:1067:4  */
  always @*
    case (n7981)
      8'b10000000: n7982 = 16'b1001101101000100;
      8'b01000000: n7982 = 16'b1000010100010110;
      8'b00100000: n7982 = 16'b0110111011100111;
      8'b00010000: n7982 = 16'b0101100010111001;
      8'b00001000: n7982 = 16'b0100001010001011;
      8'b00000100: n7982 = 16'b0010110001011101;
      8'b00000010: n7982 = 16'b0001011000101110;
      8'b00000001: n7982 = 16'b0000000000000000;
      default: n7982 = 16'bX;
    endcase
endmodule

module fixrealkcm_freq500_uid89_t0_freq500_uid92
  (input  [4:0] x,
   output [20:0] y);
  wire [20:0] y0;
  wire [20:0] y1;
  wire n7858;
  wire n7861;
  wire n7864;
  wire n7867;
  wire n7870;
  wire n7873;
  wire n7876;
  wire n7879;
  wire n7882;
  wire n7885;
  wire n7888;
  wire n7891;
  wire n7894;
  wire n7897;
  wire n7900;
  wire n7903;
  wire n7906;
  wire n7909;
  wire n7912;
  wire n7915;
  wire n7918;
  wire n7921;
  wire n7924;
  wire n7927;
  wire n7930;
  wire n7933;
  wire n7936;
  wire n7939;
  wire n7942;
  wire n7945;
  wire n7948;
  wire n7951;
  wire [31:0] n7953;
  reg [20:0] n7954;
  assign y = y1; //(module output)
  /* fppowtf32.vhdl:990:8  */
  assign y0 = n7954; // (signal)
  /* fppowtf32.vhdl:992:8  */
  assign y1 = y0; // (signal)
  /* fppowtf32.vhdl:996:31  */
  assign n7858 = x == 5'b00000;
  /* fppowtf32.vhdl:997:31  */
  assign n7861 = x == 5'b00001;
  /* fppowtf32.vhdl:998:31  */
  assign n7864 = x == 5'b00010;
  /* fppowtf32.vhdl:999:31  */
  assign n7867 = x == 5'b00011;
  /* fppowtf32.vhdl:1000:31  */
  assign n7870 = x == 5'b00100;
  /* fppowtf32.vhdl:1001:31  */
  assign n7873 = x == 5'b00101;
  /* fppowtf32.vhdl:1002:31  */
  assign n7876 = x == 5'b00110;
  /* fppowtf32.vhdl:1003:31  */
  assign n7879 = x == 5'b00111;
  /* fppowtf32.vhdl:1004:31  */
  assign n7882 = x == 5'b01000;
  /* fppowtf32.vhdl:1005:31  */
  assign n7885 = x == 5'b01001;
  /* fppowtf32.vhdl:1006:31  */
  assign n7888 = x == 5'b01010;
  /* fppowtf32.vhdl:1007:31  */
  assign n7891 = x == 5'b01011;
  /* fppowtf32.vhdl:1008:31  */
  assign n7894 = x == 5'b01100;
  /* fppowtf32.vhdl:1009:31  */
  assign n7897 = x == 5'b01101;
  /* fppowtf32.vhdl:1010:31  */
  assign n7900 = x == 5'b01110;
  /* fppowtf32.vhdl:1011:31  */
  assign n7903 = x == 5'b01111;
  /* fppowtf32.vhdl:1012:31  */
  assign n7906 = x == 5'b10000;
  /* fppowtf32.vhdl:1013:31  */
  assign n7909 = x == 5'b10001;
  /* fppowtf32.vhdl:1014:31  */
  assign n7912 = x == 5'b10010;
  /* fppowtf32.vhdl:1015:31  */
  assign n7915 = x == 5'b10011;
  /* fppowtf32.vhdl:1016:31  */
  assign n7918 = x == 5'b10100;
  /* fppowtf32.vhdl:1017:31  */
  assign n7921 = x == 5'b10101;
  /* fppowtf32.vhdl:1018:31  */
  assign n7924 = x == 5'b10110;
  /* fppowtf32.vhdl:1019:31  */
  assign n7927 = x == 5'b10111;
  /* fppowtf32.vhdl:1020:31  */
  assign n7930 = x == 5'b11000;
  /* fppowtf32.vhdl:1021:31  */
  assign n7933 = x == 5'b11001;
  /* fppowtf32.vhdl:1022:31  */
  assign n7936 = x == 5'b11010;
  /* fppowtf32.vhdl:1023:31  */
  assign n7939 = x == 5'b11011;
  /* fppowtf32.vhdl:1024:31  */
  assign n7942 = x == 5'b11100;
  /* fppowtf32.vhdl:1025:31  */
  assign n7945 = x == 5'b11101;
  /* fppowtf32.vhdl:1026:31  */
  assign n7948 = x == 5'b11110;
  /* fppowtf32.vhdl:1027:31  */
  assign n7951 = x == 5'b11111;
  assign n7953 = {n7951, n7948, n7945, n7942, n7939, n7936, n7933, n7930, n7927, n7924, n7921, n7918, n7915, n7912, n7909, n7906, n7903, n7900, n7897, n7894, n7891, n7888, n7885, n7882, n7879, n7876, n7873, n7870, n7867, n7864, n7861, n7858};
  /* fppowtf32.vhdl:995:4  */
  always @*
    case (n7953)
      32'b10000000000000000000000000000000: n7954 = 21'b101010111110011010001;
      32'b01000000000000000000000000000000: n7954 = 21'b101001100101101011111;
      32'b00100000000000000000000000000000: n7954 = 21'b101000001100111101101;
      32'b00010000000000000000000000000000: n7954 = 21'b100110110100001111011;
      32'b00001000000000000000000000000000: n7954 = 21'b100101011011100001001;
      32'b00000100000000000000000000000000: n7954 = 21'b100100000010110010110;
      32'b00000010000000000000000000000000: n7954 = 21'b100010101010000100100;
      32'b00000001000000000000000000000000: n7954 = 21'b100001010001010110010;
      32'b00000000100000000000000000000000: n7954 = 21'b011111111000101000000;
      32'b00000000010000000000000000000000: n7954 = 21'b011110011111111001110;
      32'b00000000001000000000000000000000: n7954 = 21'b011101000111001011100;
      32'b00000000000100000000000000000000: n7954 = 21'b011011101110011101010;
      32'b00000000000010000000000000000000: n7954 = 21'b011010010101101111000;
      32'b00000000000001000000000000000000: n7954 = 21'b011000111101000000110;
      32'b00000000000000100000000000000000: n7954 = 21'b010111100100010010100;
      32'b00000000000000010000000000000000: n7954 = 21'b010110001011100100001;
      32'b00000000000000001000000000000000: n7954 = 21'b010100110010110101111;
      32'b00000000000000000100000000000000: n7954 = 21'b010011011010000111101;
      32'b00000000000000000010000000000000: n7954 = 21'b010010000001011001011;
      32'b00000000000000000001000000000000: n7954 = 21'b010000101000101011001;
      32'b00000000000000000000100000000000: n7954 = 21'b001111001111111100111;
      32'b00000000000000000000010000000000: n7954 = 21'b001101110111001110101;
      32'b00000000000000000000001000000000: n7954 = 21'b001100011110100000011;
      32'b00000000000000000000000100000000: n7954 = 21'b001011000101110010001;
      32'b00000000000000000000000010000000: n7954 = 21'b001001101101000011111;
      32'b00000000000000000000000001000000: n7954 = 21'b001000010100010101101;
      32'b00000000000000000000000000100000: n7954 = 21'b000110111011100111010;
      32'b00000000000000000000000000010000: n7954 = 21'b000101100010111001000;
      32'b00000000000000000000000000001000: n7954 = 21'b000100001010001010110;
      32'b00000000000000000000000000000100: n7954 = 21'b000010110001011100100;
      32'b00000000000000000000000000000010: n7954 = 21'b000001011000101110010;
      32'b00000000000000000000000000000001: n7954 = 21'b000000000000000000000;
      default: n7954 = 21'bX;
    endcase
endmodule

module intadder_12_freq500_uid87
  (input  clk,
   input  [11:0] x,
   input  [11:0] y,
   input  cin,
   output [11:0] r);
  wire [11:0] rtmp;
  wire [11:0] x_d1;
  wire [11:0] y_d1;
  wire cin_d1;
  wire cin_d2;
  wire cin_d3;
  wire cin_d4;
  wire cin_d5;
  wire cin_d6;
  wire cin_d7;
  wire cin_d8;
  wire cin_d9;
  wire cin_d10;
  wire cin_d11;
  wire cin_d12;
  wire cin_d13;
  wire cin_d14;
  wire cin_d15;
  wire cin_d16;
  wire [11:0] n7834;
  wire [11:0] n7835;
  wire [11:0] n7836;
  reg [11:0] n7837;
  reg [11:0] n7838;
  reg n7839;
  reg n7840;
  reg n7841;
  reg n7842;
  reg n7843;
  reg n7844;
  reg n7845;
  reg n7846;
  reg n7847;
  reg n7848;
  reg n7849;
  reg n7850;
  reg n7851;
  reg n7852;
  reg n7853;
  reg n7854;
  assign r = rtmp; //(module output)
  /* fppowtf32.vhdl:4440:8  */
  assign rtmp = n7836; // (signal)
  /* fppowtf32.vhdl:4442:8  */
  assign x_d1 = n7837; // (signal)
  /* fppowtf32.vhdl:4444:8  */
  assign y_d1 = n7838; // (signal)
  /* fppowtf32.vhdl:4446:8  */
  assign cin_d1 = n7839; // (signal)
  /* fppowtf32.vhdl:4446:16  */
  assign cin_d2 = n7840; // (signal)
  /* fppowtf32.vhdl:4446:24  */
  assign cin_d3 = n7841; // (signal)
  /* fppowtf32.vhdl:4446:32  */
  assign cin_d4 = n7842; // (signal)
  /* fppowtf32.vhdl:4446:40  */
  assign cin_d5 = n7843; // (signal)
  /* fppowtf32.vhdl:4446:48  */
  assign cin_d6 = n7844; // (signal)
  /* fppowtf32.vhdl:4446:56  */
  assign cin_d7 = n7845; // (signal)
  /* fppowtf32.vhdl:4446:64  */
  assign cin_d8 = n7846; // (signal)
  /* fppowtf32.vhdl:4446:72  */
  assign cin_d9 = n7847; // (signal)
  /* fppowtf32.vhdl:4446:80  */
  assign cin_d10 = n7848; // (signal)
  /* fppowtf32.vhdl:4446:89  */
  assign cin_d11 = n7849; // (signal)
  /* fppowtf32.vhdl:4446:98  */
  assign cin_d12 = n7850; // (signal)
  /* fppowtf32.vhdl:4446:107  */
  assign cin_d13 = n7851; // (signal)
  /* fppowtf32.vhdl:4446:116  */
  assign cin_d14 = n7852; // (signal)
  /* fppowtf32.vhdl:4446:125  */
  assign cin_d15 = n7853; // (signal)
  /* fppowtf32.vhdl:4446:134  */
  assign cin_d16 = n7854; // (signal)
  /* fppowtf32.vhdl:4472:17  */
  assign n7834 = x_d1 + y_d1;
  /* fppowtf32.vhdl:4472:24  */
  assign n7835 = {11'b0, cin_d16};  //  uext
  /* fppowtf32.vhdl:4472:24  */
  assign n7836 = n7834 + n7835;
  /* fppowtf32.vhdl:4451:10  */
  always @(posedge clk)
    n7837 <= x;
  /* fppowtf32.vhdl:4451:10  */
  always @(posedge clk)
    n7838 <= y;
  /* fppowtf32.vhdl:4451:10  */
  always @(posedge clk)
    n7839 <= cin;
  /* fppowtf32.vhdl:4451:10  */
  always @(posedge clk)
    n7840 <= cin_d1;
  /* fppowtf32.vhdl:4451:10  */
  always @(posedge clk)
    n7841 <= cin_d2;
  /* fppowtf32.vhdl:4451:10  */
  always @(posedge clk)
    n7842 <= cin_d3;
  /* fppowtf32.vhdl:4451:10  */
  always @(posedge clk)
    n7843 <= cin_d4;
  /* fppowtf32.vhdl:4451:10  */
  always @(posedge clk)
    n7844 <= cin_d5;
  /* fppowtf32.vhdl:4451:10  */
  always @(posedge clk)
    n7845 <= cin_d6;
  /* fppowtf32.vhdl:4451:10  */
  always @(posedge clk)
    n7846 <= cin_d7;
  /* fppowtf32.vhdl:4451:10  */
  always @(posedge clk)
    n7847 <= cin_d8;
  /* fppowtf32.vhdl:4451:10  */
  always @(posedge clk)
    n7848 <= cin_d9;
  /* fppowtf32.vhdl:4451:10  */
  always @(posedge clk)
    n7849 <= cin_d10;
  /* fppowtf32.vhdl:4451:10  */
  always @(posedge clk)
    n7850 <= cin_d11;
  /* fppowtf32.vhdl:4451:10  */
  always @(posedge clk)
    n7851 <= cin_d12;
  /* fppowtf32.vhdl:4451:10  */
  always @(posedge clk)
    n7852 <= cin_d13;
  /* fppowtf32.vhdl:4451:10  */
  always @(posedge clk)
    n7853 <= cin_d14;
  /* fppowtf32.vhdl:4451:10  */
  always @(posedge clk)
    n7854 <= cin_d15;
endmodule

module fixrealkcm_freq500_uid77_t1_freq500_uid83
  (input  [4:0] x,
   output [6:0] y);
  wire [6:0] y0;
  wire [6:0] y1;
  wire n7714;
  wire n7717;
  wire n7720;
  wire n7723;
  wire n7726;
  wire n7729;
  wire n7732;
  wire n7735;
  wire n7738;
  wire n7741;
  wire n7744;
  wire n7747;
  wire n7750;
  wire n7753;
  wire n7756;
  wire n7759;
  wire n7762;
  wire n7765;
  wire n7768;
  wire n7771;
  wire n7774;
  wire n7777;
  wire n7780;
  wire n7783;
  wire n7786;
  wire n7789;
  wire n7792;
  wire n7795;
  wire n7798;
  wire n7801;
  wire n7804;
  wire n7807;
  wire [31:0] n7809;
  reg [6:0] n7810;
  assign y = y1; //(module output)
  /* fppowtf32.vhdl:918:8  */
  assign y0 = n7810; // (signal)
  /* fppowtf32.vhdl:920:8  */
  assign y1 = y0; // (signal)
  /* fppowtf32.vhdl:924:17  */
  assign n7714 = x == 5'b00000;
  /* fppowtf32.vhdl:925:17  */
  assign n7717 = x == 5'b00001;
  /* fppowtf32.vhdl:926:17  */
  assign n7720 = x == 5'b00010;
  /* fppowtf32.vhdl:927:17  */
  assign n7723 = x == 5'b00011;
  /* fppowtf32.vhdl:928:17  */
  assign n7726 = x == 5'b00100;
  /* fppowtf32.vhdl:929:17  */
  assign n7729 = x == 5'b00101;
  /* fppowtf32.vhdl:930:17  */
  assign n7732 = x == 5'b00110;
  /* fppowtf32.vhdl:931:17  */
  assign n7735 = x == 5'b00111;
  /* fppowtf32.vhdl:932:17  */
  assign n7738 = x == 5'b01000;
  /* fppowtf32.vhdl:933:17  */
  assign n7741 = x == 5'b01001;
  /* fppowtf32.vhdl:934:17  */
  assign n7744 = x == 5'b01010;
  /* fppowtf32.vhdl:935:17  */
  assign n7747 = x == 5'b01011;
  /* fppowtf32.vhdl:936:17  */
  assign n7750 = x == 5'b01100;
  /* fppowtf32.vhdl:937:17  */
  assign n7753 = x == 5'b01101;
  /* fppowtf32.vhdl:938:17  */
  assign n7756 = x == 5'b01110;
  /* fppowtf32.vhdl:939:17  */
  assign n7759 = x == 5'b01111;
  /* fppowtf32.vhdl:940:17  */
  assign n7762 = x == 5'b10000;
  /* fppowtf32.vhdl:941:17  */
  assign n7765 = x == 5'b10001;
  /* fppowtf32.vhdl:942:17  */
  assign n7768 = x == 5'b10010;
  /* fppowtf32.vhdl:943:17  */
  assign n7771 = x == 5'b10011;
  /* fppowtf32.vhdl:944:17  */
  assign n7774 = x == 5'b10100;
  /* fppowtf32.vhdl:945:17  */
  assign n7777 = x == 5'b10101;
  /* fppowtf32.vhdl:946:17  */
  assign n7780 = x == 5'b10110;
  /* fppowtf32.vhdl:947:17  */
  assign n7783 = x == 5'b10111;
  /* fppowtf32.vhdl:948:17  */
  assign n7786 = x == 5'b11000;
  /* fppowtf32.vhdl:949:17  */
  assign n7789 = x == 5'b11001;
  /* fppowtf32.vhdl:950:17  */
  assign n7792 = x == 5'b11010;
  /* fppowtf32.vhdl:951:17  */
  assign n7795 = x == 5'b11011;
  /* fppowtf32.vhdl:952:17  */
  assign n7798 = x == 5'b11100;
  /* fppowtf32.vhdl:953:17  */
  assign n7801 = x == 5'b11101;
  /* fppowtf32.vhdl:954:17  */
  assign n7804 = x == 5'b11110;
  /* fppowtf32.vhdl:955:17  */
  assign n7807 = x == 5'b11111;
  assign n7809 = {n7807, n7804, n7801, n7798, n7795, n7792, n7789, n7786, n7783, n7780, n7777, n7774, n7771, n7768, n7765, n7762, n7759, n7756, n7753, n7750, n7747, n7744, n7741, n7738, n7735, n7732, n7729, n7726, n7723, n7720, n7717, n7714};
  /* fppowtf32.vhdl:923:4  */
  always @*
    case (n7809)
      32'b10000000000000000000000000000000: n7810 = 7'b1011001;
      32'b01000000000000000000000000000000: n7810 = 7'b1010111;
      32'b00100000000000000000000000000000: n7810 = 7'b1010100;
      32'b00010000000000000000000000000000: n7810 = 7'b1010001;
      32'b00001000000000000000000000000000: n7810 = 7'b1001110;
      32'b00000100000000000000000000000000: n7810 = 7'b1001011;
      32'b00000010000000000000000000000000: n7810 = 7'b1001000;
      32'b00000001000000000000000000000000: n7810 = 7'b1000101;
      32'b00000000100000000000000000000000: n7810 = 7'b1000010;
      32'b00000000010000000000000000000000: n7810 = 7'b0111111;
      32'b00000000001000000000000000000000: n7810 = 7'b0111101;
      32'b00000000000100000000000000000000: n7810 = 7'b0111010;
      32'b00000000000010000000000000000000: n7810 = 7'b0110111;
      32'b00000000000001000000000000000000: n7810 = 7'b0110100;
      32'b00000000000000100000000000000000: n7810 = 7'b0110001;
      32'b00000000000000010000000000000000: n7810 = 7'b0101110;
      32'b00000000000000001000000000000000: n7810 = 7'b0101011;
      32'b00000000000000000100000000000000: n7810 = 7'b0101000;
      32'b00000000000000000010000000000000: n7810 = 7'b0100110;
      32'b00000000000000000001000000000000: n7810 = 7'b0100011;
      32'b00000000000000000000100000000000: n7810 = 7'b0100000;
      32'b00000000000000000000010000000000: n7810 = 7'b0011101;
      32'b00000000000000000000001000000000: n7810 = 7'b0011010;
      32'b00000000000000000000000100000000: n7810 = 7'b0010111;
      32'b00000000000000000000000010000000: n7810 = 7'b0010100;
      32'b00000000000000000000000001000000: n7810 = 7'b0010001;
      32'b00000000000000000000000000100000: n7810 = 7'b0001110;
      32'b00000000000000000000000000010000: n7810 = 7'b0001100;
      32'b00000000000000000000000000001000: n7810 = 7'b0001001;
      32'b00000000000000000000000000000100: n7810 = 7'b0000110;
      32'b00000000000000000000000000000010: n7810 = 7'b0000011;
      32'b00000000000000000000000000000001: n7810 = 7'b0000000;
      default: n7810 = 7'bX;
    endcase
endmodule

module fixrealkcm_freq500_uid77_t0_freq500_uid80
  (input  [4:0] x,
   output [11:0] y);
  wire [11:0] y0;
  wire [11:0] y1;
  wire n7614;
  wire n7617;
  wire n7620;
  wire n7623;
  wire n7626;
  wire n7629;
  wire n7632;
  wire n7635;
  wire n7638;
  wire n7641;
  wire n7644;
  wire n7647;
  wire n7650;
  wire n7653;
  wire n7656;
  wire n7659;
  wire n7662;
  wire n7665;
  wire n7668;
  wire n7671;
  wire n7674;
  wire n7677;
  wire n7680;
  wire n7683;
  wire n7686;
  wire n7689;
  wire n7692;
  wire n7695;
  wire n7698;
  wire n7701;
  wire n7704;
  wire n7707;
  wire [31:0] n7709;
  reg [11:0] n7710;
  assign y = y1; //(module output)
  /* fppowtf32.vhdl:846:8  */
  assign y0 = n7710; // (signal)
  /* fppowtf32.vhdl:848:8  */
  assign y1 = y0; // (signal)
  /* fppowtf32.vhdl:852:22  */
  assign n7614 = x == 5'b00000;
  /* fppowtf32.vhdl:853:22  */
  assign n7617 = x == 5'b00001;
  /* fppowtf32.vhdl:854:22  */
  assign n7620 = x == 5'b00010;
  /* fppowtf32.vhdl:855:22  */
  assign n7623 = x == 5'b00011;
  /* fppowtf32.vhdl:856:22  */
  assign n7626 = x == 5'b00100;
  /* fppowtf32.vhdl:857:22  */
  assign n7629 = x == 5'b00101;
  /* fppowtf32.vhdl:858:22  */
  assign n7632 = x == 5'b00110;
  /* fppowtf32.vhdl:859:22  */
  assign n7635 = x == 5'b00111;
  /* fppowtf32.vhdl:860:22  */
  assign n7638 = x == 5'b01000;
  /* fppowtf32.vhdl:861:22  */
  assign n7641 = x == 5'b01001;
  /* fppowtf32.vhdl:862:22  */
  assign n7644 = x == 5'b01010;
  /* fppowtf32.vhdl:863:22  */
  assign n7647 = x == 5'b01011;
  /* fppowtf32.vhdl:864:22  */
  assign n7650 = x == 5'b01100;
  /* fppowtf32.vhdl:865:22  */
  assign n7653 = x == 5'b01101;
  /* fppowtf32.vhdl:866:22  */
  assign n7656 = x == 5'b01110;
  /* fppowtf32.vhdl:867:22  */
  assign n7659 = x == 5'b01111;
  /* fppowtf32.vhdl:868:22  */
  assign n7662 = x == 5'b10000;
  /* fppowtf32.vhdl:869:22  */
  assign n7665 = x == 5'b10001;
  /* fppowtf32.vhdl:870:22  */
  assign n7668 = x == 5'b10010;
  /* fppowtf32.vhdl:871:22  */
  assign n7671 = x == 5'b10011;
  /* fppowtf32.vhdl:872:22  */
  assign n7674 = x == 5'b10100;
  /* fppowtf32.vhdl:873:22  */
  assign n7677 = x == 5'b10101;
  /* fppowtf32.vhdl:874:22  */
  assign n7680 = x == 5'b10110;
  /* fppowtf32.vhdl:875:22  */
  assign n7683 = x == 5'b10111;
  /* fppowtf32.vhdl:876:22  */
  assign n7686 = x == 5'b11000;
  /* fppowtf32.vhdl:877:22  */
  assign n7689 = x == 5'b11001;
  /* fppowtf32.vhdl:878:22  */
  assign n7692 = x == 5'b11010;
  /* fppowtf32.vhdl:879:22  */
  assign n7695 = x == 5'b11011;
  /* fppowtf32.vhdl:880:22  */
  assign n7698 = x == 5'b11100;
  /* fppowtf32.vhdl:881:22  */
  assign n7701 = x == 5'b11101;
  /* fppowtf32.vhdl:882:22  */
  assign n7704 = x == 5'b11110;
  /* fppowtf32.vhdl:883:22  */
  assign n7707 = x == 5'b11111;
  assign n7709 = {n7707, n7704, n7701, n7698, n7695, n7692, n7689, n7686, n7683, n7680, n7677, n7674, n7671, n7668, n7665, n7662, n7659, n7656, n7653, n7650, n7647, n7644, n7641, n7638, n7635, n7632, n7629, n7626, n7623, n7620, n7617, n7614};
  /* fppowtf32.vhdl:851:4  */
  always @*
    case (n7709)
      32'b10000000000000000000000000000000: n7710 = 12'b101100110110;
      32'b01000000000000000000000000000000: n7710 = 12'b101011011010;
      32'b00100000000000000000000000000000: n7710 = 12'b101001111110;
      32'b00010000000000000000000000000000: n7710 = 12'b101000100001;
      32'b00001000000000000000000000000000: n7710 = 12'b100111000101;
      32'b00000100000000000000000000000000: n7710 = 12'b100101101001;
      32'b00000010000000000000000000000000: n7710 = 12'b100100001100;
      32'b00000001000000000000000000000000: n7710 = 12'b100010110000;
      32'b00000000100000000000000000000000: n7710 = 12'b100001010100;
      32'b00000000010000000000000000000000: n7710 = 12'b011111110111;
      32'b00000000001000000000000000000000: n7710 = 12'b011110011011;
      32'b00000000000100000000000000000000: n7710 = 12'b011100111111;
      32'b00000000000010000000000000000000: n7710 = 12'b011011100010;
      32'b00000000000001000000000000000000: n7710 = 12'b011010000110;
      32'b00000000000000100000000000000000: n7710 = 12'b011000101010;
      32'b00000000000000010000000000000000: n7710 = 12'b010111001101;
      32'b00000000000000001000000000000000: n7710 = 12'b010101110001;
      32'b00000000000000000100000000000000: n7710 = 12'b010100010101;
      32'b00000000000000000010000000000000: n7710 = 12'b010010111000;
      32'b00000000000000000001000000000000: n7710 = 12'b010001011100;
      32'b00000000000000000000100000000000: n7710 = 12'b010000000000;
      32'b00000000000000000000010000000000: n7710 = 12'b001110100011;
      32'b00000000000000000000001000000000: n7710 = 12'b001101000111;
      32'b00000000000000000000000100000000: n7710 = 12'b001011101011;
      32'b00000000000000000000000010000000: n7710 = 12'b001010001110;
      32'b00000000000000000000000001000000: n7710 = 12'b001000110010;
      32'b00000000000000000000000000100000: n7710 = 12'b000111010110;
      32'b00000000000000000000000000010000: n7710 = 12'b000101111001;
      32'b00000000000000000000000000001000: n7710 = 12'b000100011101;
      32'b00000000000000000000000000000100: n7710 = 12'b000011000001;
      32'b00000000000000000000000000000010: n7710 = 12'b000001100100;
      32'b00000000000000000000000000000001: n7710 = 12'b000000001000;
      default: n7710 = 12'bX;
    endcase
endmodule

module intadder_14_freq500_uid118
  (input  clk,
   input  [13:0] x,
   input  [13:0] y,
   input  cin,
   output [13:0] r);
  wire [13:0] rtmp;
  wire [13:0] x_d1;
  wire cin_d1;
  wire cin_d2;
  wire cin_d3;
  wire cin_d4;
  wire cin_d5;
  wire cin_d6;
  wire cin_d7;
  wire cin_d8;
  wire cin_d9;
  wire cin_d10;
  wire cin_d11;
  wire cin_d12;
  wire cin_d13;
  wire cin_d14;
  wire cin_d15;
  wire cin_d16;
  wire cin_d17;
  wire cin_d18;
  wire cin_d19;
  wire [13:0] n7588;
  wire [13:0] n7589;
  wire [13:0] n7590;
  reg [13:0] n7591;
  reg n7592;
  reg n7593;
  reg n7594;
  reg n7595;
  reg n7596;
  reg n7597;
  reg n7598;
  reg n7599;
  reg n7600;
  reg n7601;
  reg n7602;
  reg n7603;
  reg n7604;
  reg n7605;
  reg n7606;
  reg n7607;
  reg n7608;
  reg n7609;
  reg n7610;
  assign r = rtmp; //(module output)
  /* fppowtf32.vhdl:5169:8  */
  assign rtmp = n7590; // (signal)
  /* fppowtf32.vhdl:5171:8  */
  assign x_d1 = n7591; // (signal)
  /* fppowtf32.vhdl:5173:8  */
  assign cin_d1 = n7592; // (signal)
  /* fppowtf32.vhdl:5173:16  */
  assign cin_d2 = n7593; // (signal)
  /* fppowtf32.vhdl:5173:24  */
  assign cin_d3 = n7594; // (signal)
  /* fppowtf32.vhdl:5173:32  */
  assign cin_d4 = n7595; // (signal)
  /* fppowtf32.vhdl:5173:40  */
  assign cin_d5 = n7596; // (signal)
  /* fppowtf32.vhdl:5173:48  */
  assign cin_d6 = n7597; // (signal)
  /* fppowtf32.vhdl:5173:56  */
  assign cin_d7 = n7598; // (signal)
  /* fppowtf32.vhdl:5173:64  */
  assign cin_d8 = n7599; // (signal)
  /* fppowtf32.vhdl:5173:72  */
  assign cin_d9 = n7600; // (signal)
  /* fppowtf32.vhdl:5173:80  */
  assign cin_d10 = n7601; // (signal)
  /* fppowtf32.vhdl:5173:89  */
  assign cin_d11 = n7602; // (signal)
  /* fppowtf32.vhdl:5173:98  */
  assign cin_d12 = n7603; // (signal)
  /* fppowtf32.vhdl:5173:107  */
  assign cin_d13 = n7604; // (signal)
  /* fppowtf32.vhdl:5173:116  */
  assign cin_d14 = n7605; // (signal)
  /* fppowtf32.vhdl:5173:125  */
  assign cin_d15 = n7606; // (signal)
  /* fppowtf32.vhdl:5173:134  */
  assign cin_d16 = n7607; // (signal)
  /* fppowtf32.vhdl:5173:143  */
  assign cin_d17 = n7608; // (signal)
  /* fppowtf32.vhdl:5173:152  */
  assign cin_d18 = n7609; // (signal)
  /* fppowtf32.vhdl:5173:161  */
  assign cin_d19 = n7610; // (signal)
  /* fppowtf32.vhdl:5201:17  */
  assign n7588 = x_d1 + y;
  /* fppowtf32.vhdl:5201:21  */
  assign n7589 = {13'b0, cin_d19};  //  uext
  /* fppowtf32.vhdl:5201:21  */
  assign n7590 = n7588 + n7589;
  /* fppowtf32.vhdl:5178:10  */
  always @(posedge clk)
    n7591 <= x;
  /* fppowtf32.vhdl:5178:10  */
  always @(posedge clk)
    n7592 <= cin;
  /* fppowtf32.vhdl:5178:10  */
  always @(posedge clk)
    n7593 <= cin_d1;
  /* fppowtf32.vhdl:5178:10  */
  always @(posedge clk)
    n7594 <= cin_d2;
  /* fppowtf32.vhdl:5178:10  */
  always @(posedge clk)
    n7595 <= cin_d3;
  /* fppowtf32.vhdl:5178:10  */
  always @(posedge clk)
    n7596 <= cin_d4;
  /* fppowtf32.vhdl:5178:10  */
  always @(posedge clk)
    n7597 <= cin_d5;
  /* fppowtf32.vhdl:5178:10  */
  always @(posedge clk)
    n7598 <= cin_d6;
  /* fppowtf32.vhdl:5178:10  */
  always @(posedge clk)
    n7599 <= cin_d7;
  /* fppowtf32.vhdl:5178:10  */
  always @(posedge clk)
    n7600 <= cin_d8;
  /* fppowtf32.vhdl:5178:10  */
  always @(posedge clk)
    n7601 <= cin_d9;
  /* fppowtf32.vhdl:5178:10  */
  always @(posedge clk)
    n7602 <= cin_d10;
  /* fppowtf32.vhdl:5178:10  */
  always @(posedge clk)
    n7603 <= cin_d11;
  /* fppowtf32.vhdl:5178:10  */
  always @(posedge clk)
    n7604 <= cin_d12;
  /* fppowtf32.vhdl:5178:10  */
  always @(posedge clk)
    n7605 <= cin_d13;
  /* fppowtf32.vhdl:5178:10  */
  always @(posedge clk)
    n7606 <= cin_d14;
  /* fppowtf32.vhdl:5178:10  */
  always @(posedge clk)
    n7607 <= cin_d15;
  /* fppowtf32.vhdl:5178:10  */
  always @(posedge clk)
    n7608 <= cin_d16;
  /* fppowtf32.vhdl:5178:10  */
  always @(posedge clk)
    n7609 <= cin_d17;
  /* fppowtf32.vhdl:5178:10  */
  always @(posedge clk)
    n7610 <= cin_d18;
endmodule

module intmultiplier_3x4_5_freq500_uid114
  (input  clk,
   input  [2:0] x,
   input  [3:0] y,
   output [4:0] r);
  wire [2:0] xx;
  wire [3:0] yy;
  wire [3:0] yy_d1;
  wire [6:0] rr;
  wire [6:0] n7558;
  wire [6:0] n7559;
  wire [6:0] n7560;
  wire [4:0] n7561;
  reg [3:0] n7562;
  assign r = n7561; //(module output)
  /* fppowtf32.vhdl:5118:12  */
  assign yy_d1 = n7562; // (signal)
  /* fppowtf32.vhdl:5120:8  */
  assign rr = n7560; // (signal)
  /* fppowtf32.vhdl:5133:12  */
  assign n7558 = {4'b0, xx};  //  uext
  /* fppowtf32.vhdl:5133:12  */
  assign n7559 = {3'b0, yy_d1};  //  uext
  /* fppowtf32.vhdl:5133:12  */
  assign n7560 = n7558 * n7559; // umul
  /* fppowtf32.vhdl:5134:28  */
  assign n7561 = rr[6:2]; // extract
  /* fppowtf32.vhdl:5125:10  */
  always @(posedge clk)
    n7562 <= yy;
endmodule

module intadder_4_freq500_uid112
  (input  clk,
   input  [3:0] x,
   input  [3:0] y,
   input  cin,
   output [3:0] r);
  wire [3:0] rtmp;
  wire [3:0] x_d1;
  wire [3:0] y_d1;
  wire [3:0] y_d2;
  wire [3:0] y_d3;
  wire [3:0] y_d4;
  wire [3:0] y_d5;
  wire [3:0] y_d6;
  wire [3:0] y_d7;
  wire [3:0] y_d8;
  wire [3:0] y_d9;
  wire [3:0] y_d10;
  wire [3:0] y_d11;
  wire [3:0] y_d12;
  wire [3:0] y_d13;
  wire [3:0] y_d14;
  wire [3:0] y_d15;
  wire [3:0] y_d16;
  wire [3:0] y_d17;
  wire [3:0] y_d18;
  wire [3:0] y_d19;
  wire cin_d1;
  wire cin_d2;
  wire cin_d3;
  wire cin_d4;
  wire cin_d5;
  wire cin_d6;
  wire cin_d7;
  wire cin_d8;
  wire cin_d9;
  wire cin_d10;
  wire cin_d11;
  wire cin_d12;
  wire cin_d13;
  wire cin_d14;
  wire cin_d15;
  wire cin_d16;
  wire cin_d17;
  wire cin_d18;
  wire cin_d19;
  wire [3:0] n7510;
  wire [3:0] n7511;
  wire [3:0] n7512;
  reg [3:0] n7513;
  reg [3:0] n7514;
  reg [3:0] n7515;
  reg [3:0] n7516;
  reg [3:0] n7517;
  reg [3:0] n7518;
  reg [3:0] n7519;
  reg [3:0] n7520;
  reg [3:0] n7521;
  reg [3:0] n7522;
  reg [3:0] n7523;
  reg [3:0] n7524;
  reg [3:0] n7525;
  reg [3:0] n7526;
  reg [3:0] n7527;
  reg [3:0] n7528;
  reg [3:0] n7529;
  reg [3:0] n7530;
  reg [3:0] n7531;
  reg [3:0] n7532;
  reg n7533;
  reg n7534;
  reg n7535;
  reg n7536;
  reg n7537;
  reg n7538;
  reg n7539;
  reg n7540;
  reg n7541;
  reg n7542;
  reg n7543;
  reg n7544;
  reg n7545;
  reg n7546;
  reg n7547;
  reg n7548;
  reg n7549;
  reg n7550;
  reg n7551;
  assign r = rtmp; //(module output)
  /* fppowtf32.vhdl:5025:8  */
  assign rtmp = n7512; // (signal)
  /* fppowtf32.vhdl:5027:8  */
  assign x_d1 = n7513; // (signal)
  /* fppowtf32.vhdl:5029:8  */
  assign y_d1 = n7514; // (signal)
  /* fppowtf32.vhdl:5029:14  */
  assign y_d2 = n7515; // (signal)
  /* fppowtf32.vhdl:5029:20  */
  assign y_d3 = n7516; // (signal)
  /* fppowtf32.vhdl:5029:26  */
  assign y_d4 = n7517; // (signal)
  /* fppowtf32.vhdl:5029:32  */
  assign y_d5 = n7518; // (signal)
  /* fppowtf32.vhdl:5029:38  */
  assign y_d6 = n7519; // (signal)
  /* fppowtf32.vhdl:5029:44  */
  assign y_d7 = n7520; // (signal)
  /* fppowtf32.vhdl:5029:50  */
  assign y_d8 = n7521; // (signal)
  /* fppowtf32.vhdl:5029:56  */
  assign y_d9 = n7522; // (signal)
  /* fppowtf32.vhdl:5029:62  */
  assign y_d10 = n7523; // (signal)
  /* fppowtf32.vhdl:5029:69  */
  assign y_d11 = n7524; // (signal)
  /* fppowtf32.vhdl:5029:76  */
  assign y_d12 = n7525; // (signal)
  /* fppowtf32.vhdl:5029:83  */
  assign y_d13 = n7526; // (signal)
  /* fppowtf32.vhdl:5029:90  */
  assign y_d14 = n7527; // (signal)
  /* fppowtf32.vhdl:5029:97  */
  assign y_d15 = n7528; // (signal)
  /* fppowtf32.vhdl:5029:104  */
  assign y_d16 = n7529; // (signal)
  /* fppowtf32.vhdl:5029:111  */
  assign y_d17 = n7530; // (signal)
  /* fppowtf32.vhdl:5029:118  */
  assign y_d18 = n7531; // (signal)
  /* fppowtf32.vhdl:5029:125  */
  assign y_d19 = n7532; // (signal)
  /* fppowtf32.vhdl:5031:8  */
  assign cin_d1 = n7533; // (signal)
  /* fppowtf32.vhdl:5031:16  */
  assign cin_d2 = n7534; // (signal)
  /* fppowtf32.vhdl:5031:24  */
  assign cin_d3 = n7535; // (signal)
  /* fppowtf32.vhdl:5031:32  */
  assign cin_d4 = n7536; // (signal)
  /* fppowtf32.vhdl:5031:40  */
  assign cin_d5 = n7537; // (signal)
  /* fppowtf32.vhdl:5031:48  */
  assign cin_d6 = n7538; // (signal)
  /* fppowtf32.vhdl:5031:56  */
  assign cin_d7 = n7539; // (signal)
  /* fppowtf32.vhdl:5031:64  */
  assign cin_d8 = n7540; // (signal)
  /* fppowtf32.vhdl:5031:72  */
  assign cin_d9 = n7541; // (signal)
  /* fppowtf32.vhdl:5031:80  */
  assign cin_d10 = n7542; // (signal)
  /* fppowtf32.vhdl:5031:89  */
  assign cin_d11 = n7543; // (signal)
  /* fppowtf32.vhdl:5031:98  */
  assign cin_d12 = n7544; // (signal)
  /* fppowtf32.vhdl:5031:107  */
  assign cin_d13 = n7545; // (signal)
  /* fppowtf32.vhdl:5031:116  */
  assign cin_d14 = n7546; // (signal)
  /* fppowtf32.vhdl:5031:125  */
  assign cin_d15 = n7547; // (signal)
  /* fppowtf32.vhdl:5031:134  */
  assign cin_d16 = n7548; // (signal)
  /* fppowtf32.vhdl:5031:143  */
  assign cin_d17 = n7549; // (signal)
  /* fppowtf32.vhdl:5031:152  */
  assign cin_d18 = n7550; // (signal)
  /* fppowtf32.vhdl:5031:161  */
  assign cin_d19 = n7551; // (signal)
  /* fppowtf32.vhdl:5078:17  */
  assign n7510 = x_d1 + y_d19;
  /* fppowtf32.vhdl:5078:25  */
  assign n7511 = {3'b0, cin_d19};  //  uext
  /* fppowtf32.vhdl:5078:25  */
  assign n7512 = n7510 + n7511;
  /* fppowtf32.vhdl:5036:10  */
  always @(posedge clk)
    n7513 <= x;
  /* fppowtf32.vhdl:5036:10  */
  always @(posedge clk)
    n7514 <= y;
  /* fppowtf32.vhdl:5036:10  */
  always @(posedge clk)
    n7515 <= y_d1;
  /* fppowtf32.vhdl:5036:10  */
  always @(posedge clk)
    n7516 <= y_d2;
  /* fppowtf32.vhdl:5036:10  */
  always @(posedge clk)
    n7517 <= y_d3;
  /* fppowtf32.vhdl:5036:10  */
  always @(posedge clk)
    n7518 <= y_d4;
  /* fppowtf32.vhdl:5036:10  */
  always @(posedge clk)
    n7519 <= y_d5;
  /* fppowtf32.vhdl:5036:10  */
  always @(posedge clk)
    n7520 <= y_d6;
  /* fppowtf32.vhdl:5036:10  */
  always @(posedge clk)
    n7521 <= y_d7;
  /* fppowtf32.vhdl:5036:10  */
  always @(posedge clk)
    n7522 <= y_d8;
  /* fppowtf32.vhdl:5036:10  */
  always @(posedge clk)
    n7523 <= y_d9;
  /* fppowtf32.vhdl:5036:10  */
  always @(posedge clk)
    n7524 <= y_d10;
  /* fppowtf32.vhdl:5036:10  */
  always @(posedge clk)
    n7525 <= y_d11;
  /* fppowtf32.vhdl:5036:10  */
  always @(posedge clk)
    n7526 <= y_d12;
  /* fppowtf32.vhdl:5036:10  */
  always @(posedge clk)
    n7527 <= y_d13;
  /* fppowtf32.vhdl:5036:10  */
  always @(posedge clk)
    n7528 <= y_d14;
  /* fppowtf32.vhdl:5036:10  */
  always @(posedge clk)
    n7529 <= y_d15;
  /* fppowtf32.vhdl:5036:10  */
  always @(posedge clk)
    n7530 <= y_d16;
  /* fppowtf32.vhdl:5036:10  */
  always @(posedge clk)
    n7531 <= y_d17;
  /* fppowtf32.vhdl:5036:10  */
  always @(posedge clk)
    n7532 <= y_d18;
  /* fppowtf32.vhdl:5036:10  */
  always @(posedge clk)
    n7533 <= cin;
  /* fppowtf32.vhdl:5036:10  */
  always @(posedge clk)
    n7534 <= cin_d1;
  /* fppowtf32.vhdl:5036:10  */
  always @(posedge clk)
    n7535 <= cin_d2;
  /* fppowtf32.vhdl:5036:10  */
  always @(posedge clk)
    n7536 <= cin_d3;
  /* fppowtf32.vhdl:5036:10  */
  always @(posedge clk)
    n7537 <= cin_d4;
  /* fppowtf32.vhdl:5036:10  */
  always @(posedge clk)
    n7538 <= cin_d5;
  /* fppowtf32.vhdl:5036:10  */
  always @(posedge clk)
    n7539 <= cin_d6;
  /* fppowtf32.vhdl:5036:10  */
  always @(posedge clk)
    n7540 <= cin_d7;
  /* fppowtf32.vhdl:5036:10  */
  always @(posedge clk)
    n7541 <= cin_d8;
  /* fppowtf32.vhdl:5036:10  */
  always @(posedge clk)
    n7542 <= cin_d9;
  /* fppowtf32.vhdl:5036:10  */
  always @(posedge clk)
    n7543 <= cin_d10;
  /* fppowtf32.vhdl:5036:10  */
  always @(posedge clk)
    n7544 <= cin_d11;
  /* fppowtf32.vhdl:5036:10  */
  always @(posedge clk)
    n7545 <= cin_d12;
  /* fppowtf32.vhdl:5036:10  */
  always @(posedge clk)
    n7546 <= cin_d13;
  /* fppowtf32.vhdl:5036:10  */
  always @(posedge clk)
    n7547 <= cin_d14;
  /* fppowtf32.vhdl:5036:10  */
  always @(posedge clk)
    n7548 <= cin_d15;
  /* fppowtf32.vhdl:5036:10  */
  always @(posedge clk)
    n7549 <= cin_d16;
  /* fppowtf32.vhdl:5036:10  */
  always @(posedge clk)
    n7550 <= cin_d17;
  /* fppowtf32.vhdl:5036:10  */
  always @(posedge clk)
    n7551 <= cin_d18;
endmodule

module fixfunctionbytable_freq500_uid107
  (input  [2:0] x,
   output [2:0] y);
  wire [2:0] y0;
  wire [2:0] y1;
  wire n7441;
  wire n7444;
  wire n7447;
  wire n7450;
  wire n7453;
  wire n7456;
  wire n7459;
  wire n7462;
  wire [7:0] n7464;
  reg [2:0] n7465;
  assign y = y1; //(module output)
  /* fppowtf32.vhdl:2178:8  */
  assign y0 = n7465; // (signal)
  /* fppowtf32.vhdl:2180:8  */
  assign y1 = y0; // (signal)
  /* fppowtf32.vhdl:2184:13  */
  assign n7441 = x == 3'b000;
  /* fppowtf32.vhdl:2185:13  */
  assign n7444 = x == 3'b001;
  /* fppowtf32.vhdl:2186:13  */
  assign n7447 = x == 3'b010;
  /* fppowtf32.vhdl:2187:13  */
  assign n7450 = x == 3'b011;
  /* fppowtf32.vhdl:2188:13  */
  assign n7453 = x == 3'b100;
  /* fppowtf32.vhdl:2189:13  */
  assign n7456 = x == 3'b101;
  /* fppowtf32.vhdl:2190:13  */
  assign n7459 = x == 3'b110;
  /* fppowtf32.vhdl:2191:13  */
  assign n7462 = x == 3'b111;
  assign n7464 = {n7462, n7459, n7456, n7453, n7450, n7447, n7444, n7441};
  /* fppowtf32.vhdl:2183:4  */
  always @*
    case (n7464)
      8'b10000000: n7465 = 3'b111;
      8'b01000000: n7465 = 3'b110;
      8'b00100000: n7465 = 3'b101;
      8'b00010000: n7465 = 3'b100;
      8'b00001000: n7465 = 3'b011;
      8'b00000100: n7465 = 3'b010;
      8'b00000010: n7465 = 3'b001;
      8'b00000001: n7465 = 3'b000;
      default: n7465 = 3'bX;
    endcase
endmodule

module fixfunctionbytable_freq500_uid104
  (input  [9:0] x,
   output [13:0] y);
  wire [13:0] y0;
  wire [13:0] y1;
  wire n4365;
  wire n4368;
  wire n4371;
  wire n4374;
  wire n4377;
  wire n4380;
  wire n4383;
  wire n4386;
  wire n4389;
  wire n4392;
  wire n4395;
  wire n4398;
  wire n4401;
  wire n4404;
  wire n4407;
  wire n4410;
  wire n4413;
  wire n4416;
  wire n4419;
  wire n4422;
  wire n4425;
  wire n4428;
  wire n4431;
  wire n4434;
  wire n4437;
  wire n4440;
  wire n4443;
  wire n4446;
  wire n4449;
  wire n4452;
  wire n4455;
  wire n4458;
  wire n4461;
  wire n4464;
  wire n4467;
  wire n4470;
  wire n4473;
  wire n4476;
  wire n4479;
  wire n4482;
  wire n4485;
  wire n4488;
  wire n4491;
  wire n4494;
  wire n4497;
  wire n4500;
  wire n4503;
  wire n4506;
  wire n4509;
  wire n4512;
  wire n4515;
  wire n4518;
  wire n4521;
  wire n4524;
  wire n4527;
  wire n4530;
  wire n4533;
  wire n4536;
  wire n4539;
  wire n4542;
  wire n4545;
  wire n4548;
  wire n4551;
  wire n4554;
  wire n4557;
  wire n4560;
  wire n4563;
  wire n4566;
  wire n4569;
  wire n4572;
  wire n4575;
  wire n4578;
  wire n4581;
  wire n4584;
  wire n4587;
  wire n4590;
  wire n4593;
  wire n4596;
  wire n4599;
  wire n4602;
  wire n4605;
  wire n4608;
  wire n4611;
  wire n4614;
  wire n4617;
  wire n4620;
  wire n4623;
  wire n4626;
  wire n4629;
  wire n4632;
  wire n4635;
  wire n4638;
  wire n4641;
  wire n4644;
  wire n4647;
  wire n4650;
  wire n4653;
  wire n4656;
  wire n4659;
  wire n4662;
  wire n4665;
  wire n4668;
  wire n4671;
  wire n4674;
  wire n4677;
  wire n4680;
  wire n4683;
  wire n4686;
  wire n4689;
  wire n4692;
  wire n4695;
  wire n4698;
  wire n4701;
  wire n4704;
  wire n4707;
  wire n4710;
  wire n4713;
  wire n4716;
  wire n4719;
  wire n4722;
  wire n4725;
  wire n4728;
  wire n4731;
  wire n4734;
  wire n4737;
  wire n4740;
  wire n4743;
  wire n4746;
  wire n4749;
  wire n4752;
  wire n4755;
  wire n4758;
  wire n4761;
  wire n4764;
  wire n4767;
  wire n4770;
  wire n4773;
  wire n4776;
  wire n4779;
  wire n4782;
  wire n4785;
  wire n4788;
  wire n4791;
  wire n4794;
  wire n4797;
  wire n4800;
  wire n4803;
  wire n4806;
  wire n4809;
  wire n4812;
  wire n4815;
  wire n4818;
  wire n4821;
  wire n4824;
  wire n4827;
  wire n4830;
  wire n4833;
  wire n4836;
  wire n4839;
  wire n4842;
  wire n4845;
  wire n4848;
  wire n4851;
  wire n4854;
  wire n4857;
  wire n4860;
  wire n4863;
  wire n4866;
  wire n4869;
  wire n4872;
  wire n4875;
  wire n4878;
  wire n4881;
  wire n4884;
  wire n4887;
  wire n4890;
  wire n4893;
  wire n4896;
  wire n4899;
  wire n4902;
  wire n4905;
  wire n4908;
  wire n4911;
  wire n4914;
  wire n4917;
  wire n4920;
  wire n4923;
  wire n4926;
  wire n4929;
  wire n4932;
  wire n4935;
  wire n4938;
  wire n4941;
  wire n4944;
  wire n4947;
  wire n4950;
  wire n4953;
  wire n4956;
  wire n4959;
  wire n4962;
  wire n4965;
  wire n4968;
  wire n4971;
  wire n4974;
  wire n4977;
  wire n4980;
  wire n4983;
  wire n4986;
  wire n4989;
  wire n4992;
  wire n4995;
  wire n4998;
  wire n5001;
  wire n5004;
  wire n5007;
  wire n5010;
  wire n5013;
  wire n5016;
  wire n5019;
  wire n5022;
  wire n5025;
  wire n5028;
  wire n5031;
  wire n5034;
  wire n5037;
  wire n5040;
  wire n5043;
  wire n5046;
  wire n5049;
  wire n5052;
  wire n5055;
  wire n5058;
  wire n5061;
  wire n5064;
  wire n5067;
  wire n5070;
  wire n5073;
  wire n5076;
  wire n5079;
  wire n5082;
  wire n5085;
  wire n5088;
  wire n5091;
  wire n5094;
  wire n5097;
  wire n5100;
  wire n5103;
  wire n5106;
  wire n5109;
  wire n5112;
  wire n5115;
  wire n5118;
  wire n5121;
  wire n5124;
  wire n5127;
  wire n5130;
  wire n5133;
  wire n5136;
  wire n5139;
  wire n5142;
  wire n5145;
  wire n5148;
  wire n5151;
  wire n5154;
  wire n5157;
  wire n5160;
  wire n5163;
  wire n5166;
  wire n5169;
  wire n5172;
  wire n5175;
  wire n5178;
  wire n5181;
  wire n5184;
  wire n5187;
  wire n5190;
  wire n5193;
  wire n5196;
  wire n5199;
  wire n5202;
  wire n5205;
  wire n5208;
  wire n5211;
  wire n5214;
  wire n5217;
  wire n5220;
  wire n5223;
  wire n5226;
  wire n5229;
  wire n5232;
  wire n5235;
  wire n5238;
  wire n5241;
  wire n5244;
  wire n5247;
  wire n5250;
  wire n5253;
  wire n5256;
  wire n5259;
  wire n5262;
  wire n5265;
  wire n5268;
  wire n5271;
  wire n5274;
  wire n5277;
  wire n5280;
  wire n5283;
  wire n5286;
  wire n5289;
  wire n5292;
  wire n5295;
  wire n5298;
  wire n5301;
  wire n5304;
  wire n5307;
  wire n5310;
  wire n5313;
  wire n5316;
  wire n5319;
  wire n5322;
  wire n5325;
  wire n5328;
  wire n5331;
  wire n5334;
  wire n5337;
  wire n5340;
  wire n5343;
  wire n5346;
  wire n5349;
  wire n5352;
  wire n5355;
  wire n5358;
  wire n5361;
  wire n5364;
  wire n5367;
  wire n5370;
  wire n5373;
  wire n5376;
  wire n5379;
  wire n5382;
  wire n5385;
  wire n5388;
  wire n5391;
  wire n5394;
  wire n5397;
  wire n5400;
  wire n5403;
  wire n5406;
  wire n5409;
  wire n5412;
  wire n5415;
  wire n5418;
  wire n5421;
  wire n5424;
  wire n5427;
  wire n5430;
  wire n5433;
  wire n5436;
  wire n5439;
  wire n5442;
  wire n5445;
  wire n5448;
  wire n5451;
  wire n5454;
  wire n5457;
  wire n5460;
  wire n5463;
  wire n5466;
  wire n5469;
  wire n5472;
  wire n5475;
  wire n5478;
  wire n5481;
  wire n5484;
  wire n5487;
  wire n5490;
  wire n5493;
  wire n5496;
  wire n5499;
  wire n5502;
  wire n5505;
  wire n5508;
  wire n5511;
  wire n5514;
  wire n5517;
  wire n5520;
  wire n5523;
  wire n5526;
  wire n5529;
  wire n5532;
  wire n5535;
  wire n5538;
  wire n5541;
  wire n5544;
  wire n5547;
  wire n5550;
  wire n5553;
  wire n5556;
  wire n5559;
  wire n5562;
  wire n5565;
  wire n5568;
  wire n5571;
  wire n5574;
  wire n5577;
  wire n5580;
  wire n5583;
  wire n5586;
  wire n5589;
  wire n5592;
  wire n5595;
  wire n5598;
  wire n5601;
  wire n5604;
  wire n5607;
  wire n5610;
  wire n5613;
  wire n5616;
  wire n5619;
  wire n5622;
  wire n5625;
  wire n5628;
  wire n5631;
  wire n5634;
  wire n5637;
  wire n5640;
  wire n5643;
  wire n5646;
  wire n5649;
  wire n5652;
  wire n5655;
  wire n5658;
  wire n5661;
  wire n5664;
  wire n5667;
  wire n5670;
  wire n5673;
  wire n5676;
  wire n5679;
  wire n5682;
  wire n5685;
  wire n5688;
  wire n5691;
  wire n5694;
  wire n5697;
  wire n5700;
  wire n5703;
  wire n5706;
  wire n5709;
  wire n5712;
  wire n5715;
  wire n5718;
  wire n5721;
  wire n5724;
  wire n5727;
  wire n5730;
  wire n5733;
  wire n5736;
  wire n5739;
  wire n5742;
  wire n5745;
  wire n5748;
  wire n5751;
  wire n5754;
  wire n5757;
  wire n5760;
  wire n5763;
  wire n5766;
  wire n5769;
  wire n5772;
  wire n5775;
  wire n5778;
  wire n5781;
  wire n5784;
  wire n5787;
  wire n5790;
  wire n5793;
  wire n5796;
  wire n5799;
  wire n5802;
  wire n5805;
  wire n5808;
  wire n5811;
  wire n5814;
  wire n5817;
  wire n5820;
  wire n5823;
  wire n5826;
  wire n5829;
  wire n5832;
  wire n5835;
  wire n5838;
  wire n5841;
  wire n5844;
  wire n5847;
  wire n5850;
  wire n5853;
  wire n5856;
  wire n5859;
  wire n5862;
  wire n5865;
  wire n5868;
  wire n5871;
  wire n5874;
  wire n5877;
  wire n5880;
  wire n5883;
  wire n5886;
  wire n5889;
  wire n5892;
  wire n5895;
  wire n5898;
  wire n5901;
  wire n5904;
  wire n5907;
  wire n5910;
  wire n5913;
  wire n5916;
  wire n5919;
  wire n5922;
  wire n5925;
  wire n5928;
  wire n5931;
  wire n5934;
  wire n5937;
  wire n5940;
  wire n5943;
  wire n5946;
  wire n5949;
  wire n5952;
  wire n5955;
  wire n5958;
  wire n5961;
  wire n5964;
  wire n5967;
  wire n5970;
  wire n5973;
  wire n5976;
  wire n5979;
  wire n5982;
  wire n5985;
  wire n5988;
  wire n5991;
  wire n5994;
  wire n5997;
  wire n6000;
  wire n6003;
  wire n6006;
  wire n6009;
  wire n6012;
  wire n6015;
  wire n6018;
  wire n6021;
  wire n6024;
  wire n6027;
  wire n6030;
  wire n6033;
  wire n6036;
  wire n6039;
  wire n6042;
  wire n6045;
  wire n6048;
  wire n6051;
  wire n6054;
  wire n6057;
  wire n6060;
  wire n6063;
  wire n6066;
  wire n6069;
  wire n6072;
  wire n6075;
  wire n6078;
  wire n6081;
  wire n6084;
  wire n6087;
  wire n6090;
  wire n6093;
  wire n6096;
  wire n6099;
  wire n6102;
  wire n6105;
  wire n6108;
  wire n6111;
  wire n6114;
  wire n6117;
  wire n6120;
  wire n6123;
  wire n6126;
  wire n6129;
  wire n6132;
  wire n6135;
  wire n6138;
  wire n6141;
  wire n6144;
  wire n6147;
  wire n6150;
  wire n6153;
  wire n6156;
  wire n6159;
  wire n6162;
  wire n6165;
  wire n6168;
  wire n6171;
  wire n6174;
  wire n6177;
  wire n6180;
  wire n6183;
  wire n6186;
  wire n6189;
  wire n6192;
  wire n6195;
  wire n6198;
  wire n6201;
  wire n6204;
  wire n6207;
  wire n6210;
  wire n6213;
  wire n6216;
  wire n6219;
  wire n6222;
  wire n6225;
  wire n6228;
  wire n6231;
  wire n6234;
  wire n6237;
  wire n6240;
  wire n6243;
  wire n6246;
  wire n6249;
  wire n6252;
  wire n6255;
  wire n6258;
  wire n6261;
  wire n6264;
  wire n6267;
  wire n6270;
  wire n6273;
  wire n6276;
  wire n6279;
  wire n6282;
  wire n6285;
  wire n6288;
  wire n6291;
  wire n6294;
  wire n6297;
  wire n6300;
  wire n6303;
  wire n6306;
  wire n6309;
  wire n6312;
  wire n6315;
  wire n6318;
  wire n6321;
  wire n6324;
  wire n6327;
  wire n6330;
  wire n6333;
  wire n6336;
  wire n6339;
  wire n6342;
  wire n6345;
  wire n6348;
  wire n6351;
  wire n6354;
  wire n6357;
  wire n6360;
  wire n6363;
  wire n6366;
  wire n6369;
  wire n6372;
  wire n6375;
  wire n6378;
  wire n6381;
  wire n6384;
  wire n6387;
  wire n6390;
  wire n6393;
  wire n6396;
  wire n6399;
  wire n6402;
  wire n6405;
  wire n6408;
  wire n6411;
  wire n6414;
  wire n6417;
  wire n6420;
  wire n6423;
  wire n6426;
  wire n6429;
  wire n6432;
  wire n6435;
  wire n6438;
  wire n6441;
  wire n6444;
  wire n6447;
  wire n6450;
  wire n6453;
  wire n6456;
  wire n6459;
  wire n6462;
  wire n6465;
  wire n6468;
  wire n6471;
  wire n6474;
  wire n6477;
  wire n6480;
  wire n6483;
  wire n6486;
  wire n6489;
  wire n6492;
  wire n6495;
  wire n6498;
  wire n6501;
  wire n6504;
  wire n6507;
  wire n6510;
  wire n6513;
  wire n6516;
  wire n6519;
  wire n6522;
  wire n6525;
  wire n6528;
  wire n6531;
  wire n6534;
  wire n6537;
  wire n6540;
  wire n6543;
  wire n6546;
  wire n6549;
  wire n6552;
  wire n6555;
  wire n6558;
  wire n6561;
  wire n6564;
  wire n6567;
  wire n6570;
  wire n6573;
  wire n6576;
  wire n6579;
  wire n6582;
  wire n6585;
  wire n6588;
  wire n6591;
  wire n6594;
  wire n6597;
  wire n6600;
  wire n6603;
  wire n6606;
  wire n6609;
  wire n6612;
  wire n6615;
  wire n6618;
  wire n6621;
  wire n6624;
  wire n6627;
  wire n6630;
  wire n6633;
  wire n6636;
  wire n6639;
  wire n6642;
  wire n6645;
  wire n6648;
  wire n6651;
  wire n6654;
  wire n6657;
  wire n6660;
  wire n6663;
  wire n6666;
  wire n6669;
  wire n6672;
  wire n6675;
  wire n6678;
  wire n6681;
  wire n6684;
  wire n6687;
  wire n6690;
  wire n6693;
  wire n6696;
  wire n6699;
  wire n6702;
  wire n6705;
  wire n6708;
  wire n6711;
  wire n6714;
  wire n6717;
  wire n6720;
  wire n6723;
  wire n6726;
  wire n6729;
  wire n6732;
  wire n6735;
  wire n6738;
  wire n6741;
  wire n6744;
  wire n6747;
  wire n6750;
  wire n6753;
  wire n6756;
  wire n6759;
  wire n6762;
  wire n6765;
  wire n6768;
  wire n6771;
  wire n6774;
  wire n6777;
  wire n6780;
  wire n6783;
  wire n6786;
  wire n6789;
  wire n6792;
  wire n6795;
  wire n6798;
  wire n6801;
  wire n6804;
  wire n6807;
  wire n6810;
  wire n6813;
  wire n6816;
  wire n6819;
  wire n6822;
  wire n6825;
  wire n6828;
  wire n6831;
  wire n6834;
  wire n6837;
  wire n6840;
  wire n6843;
  wire n6846;
  wire n6849;
  wire n6852;
  wire n6855;
  wire n6858;
  wire n6861;
  wire n6864;
  wire n6867;
  wire n6870;
  wire n6873;
  wire n6876;
  wire n6879;
  wire n6882;
  wire n6885;
  wire n6888;
  wire n6891;
  wire n6894;
  wire n6897;
  wire n6900;
  wire n6903;
  wire n6906;
  wire n6909;
  wire n6912;
  wire n6915;
  wire n6918;
  wire n6921;
  wire n6924;
  wire n6927;
  wire n6930;
  wire n6933;
  wire n6936;
  wire n6939;
  wire n6942;
  wire n6945;
  wire n6948;
  wire n6951;
  wire n6954;
  wire n6957;
  wire n6960;
  wire n6963;
  wire n6966;
  wire n6969;
  wire n6972;
  wire n6975;
  wire n6978;
  wire n6981;
  wire n6984;
  wire n6987;
  wire n6990;
  wire n6993;
  wire n6996;
  wire n6999;
  wire n7002;
  wire n7005;
  wire n7008;
  wire n7011;
  wire n7014;
  wire n7017;
  wire n7020;
  wire n7023;
  wire n7026;
  wire n7029;
  wire n7032;
  wire n7035;
  wire n7038;
  wire n7041;
  wire n7044;
  wire n7047;
  wire n7050;
  wire n7053;
  wire n7056;
  wire n7059;
  wire n7062;
  wire n7065;
  wire n7068;
  wire n7071;
  wire n7074;
  wire n7077;
  wire n7080;
  wire n7083;
  wire n7086;
  wire n7089;
  wire n7092;
  wire n7095;
  wire n7098;
  wire n7101;
  wire n7104;
  wire n7107;
  wire n7110;
  wire n7113;
  wire n7116;
  wire n7119;
  wire n7122;
  wire n7125;
  wire n7128;
  wire n7131;
  wire n7134;
  wire n7137;
  wire n7140;
  wire n7143;
  wire n7146;
  wire n7149;
  wire n7152;
  wire n7155;
  wire n7158;
  wire n7161;
  wire n7164;
  wire n7167;
  wire n7170;
  wire n7173;
  wire n7176;
  wire n7179;
  wire n7182;
  wire n7185;
  wire n7188;
  wire n7191;
  wire n7194;
  wire n7197;
  wire n7200;
  wire n7203;
  wire n7206;
  wire n7209;
  wire n7212;
  wire n7215;
  wire n7218;
  wire n7221;
  wire n7224;
  wire n7227;
  wire n7230;
  wire n7233;
  wire n7236;
  wire n7239;
  wire n7242;
  wire n7245;
  wire n7248;
  wire n7251;
  wire n7254;
  wire n7257;
  wire n7260;
  wire n7263;
  wire n7266;
  wire n7269;
  wire n7272;
  wire n7275;
  wire n7278;
  wire n7281;
  wire n7284;
  wire n7287;
  wire n7290;
  wire n7293;
  wire n7296;
  wire n7299;
  wire n7302;
  wire n7305;
  wire n7308;
  wire n7311;
  wire n7314;
  wire n7317;
  wire n7320;
  wire n7323;
  wire n7326;
  wire n7329;
  wire n7332;
  wire n7335;
  wire n7338;
  wire n7341;
  wire n7344;
  wire n7347;
  wire n7350;
  wire n7353;
  wire n7356;
  wire n7359;
  wire n7362;
  wire n7365;
  wire n7368;
  wire n7371;
  wire n7374;
  wire n7377;
  wire n7380;
  wire n7383;
  wire n7386;
  wire n7389;
  wire n7392;
  wire n7395;
  wire n7398;
  wire n7401;
  wire n7404;
  wire n7407;
  wire n7410;
  wire n7413;
  wire n7416;
  wire n7419;
  wire n7422;
  wire n7425;
  wire n7428;
  wire n7431;
  wire n7434;
  wire [1023:0] n7436;
  reg [13:0] n7437;
  assign y = y1; //(module output)
  /* fppowtf32.vhdl:1112:8  */
  assign y0 = n7437; // (signal)
  /* fppowtf32.vhdl:1114:8  */
  assign y1 = y0; // (signal)
  /* fppowtf32.vhdl:1118:24  */
  assign n4365 = x == 10'b0000000000;
  /* fppowtf32.vhdl:1119:24  */
  assign n4368 = x == 10'b0000000001;
  /* fppowtf32.vhdl:1120:24  */
  assign n4371 = x == 10'b0000000010;
  /* fppowtf32.vhdl:1121:24  */
  assign n4374 = x == 10'b0000000011;
  /* fppowtf32.vhdl:1122:24  */
  assign n4377 = x == 10'b0000000100;
  /* fppowtf32.vhdl:1123:24  */
  assign n4380 = x == 10'b0000000101;
  /* fppowtf32.vhdl:1124:24  */
  assign n4383 = x == 10'b0000000110;
  /* fppowtf32.vhdl:1125:24  */
  assign n4386 = x == 10'b0000000111;
  /* fppowtf32.vhdl:1126:24  */
  assign n4389 = x == 10'b0000001000;
  /* fppowtf32.vhdl:1127:24  */
  assign n4392 = x == 10'b0000001001;
  /* fppowtf32.vhdl:1128:24  */
  assign n4395 = x == 10'b0000001010;
  /* fppowtf32.vhdl:1129:24  */
  assign n4398 = x == 10'b0000001011;
  /* fppowtf32.vhdl:1130:24  */
  assign n4401 = x == 10'b0000001100;
  /* fppowtf32.vhdl:1131:24  */
  assign n4404 = x == 10'b0000001101;
  /* fppowtf32.vhdl:1132:24  */
  assign n4407 = x == 10'b0000001110;
  /* fppowtf32.vhdl:1133:24  */
  assign n4410 = x == 10'b0000001111;
  /* fppowtf32.vhdl:1134:24  */
  assign n4413 = x == 10'b0000010000;
  /* fppowtf32.vhdl:1135:24  */
  assign n4416 = x == 10'b0000010001;
  /* fppowtf32.vhdl:1136:24  */
  assign n4419 = x == 10'b0000010010;
  /* fppowtf32.vhdl:1137:24  */
  assign n4422 = x == 10'b0000010011;
  /* fppowtf32.vhdl:1138:24  */
  assign n4425 = x == 10'b0000010100;
  /* fppowtf32.vhdl:1139:24  */
  assign n4428 = x == 10'b0000010101;
  /* fppowtf32.vhdl:1140:24  */
  assign n4431 = x == 10'b0000010110;
  /* fppowtf32.vhdl:1141:24  */
  assign n4434 = x == 10'b0000010111;
  /* fppowtf32.vhdl:1142:24  */
  assign n4437 = x == 10'b0000011000;
  /* fppowtf32.vhdl:1143:24  */
  assign n4440 = x == 10'b0000011001;
  /* fppowtf32.vhdl:1144:24  */
  assign n4443 = x == 10'b0000011010;
  /* fppowtf32.vhdl:1145:24  */
  assign n4446 = x == 10'b0000011011;
  /* fppowtf32.vhdl:1146:24  */
  assign n4449 = x == 10'b0000011100;
  /* fppowtf32.vhdl:1147:24  */
  assign n4452 = x == 10'b0000011101;
  /* fppowtf32.vhdl:1148:24  */
  assign n4455 = x == 10'b0000011110;
  /* fppowtf32.vhdl:1149:24  */
  assign n4458 = x == 10'b0000011111;
  /* fppowtf32.vhdl:1150:24  */
  assign n4461 = x == 10'b0000100000;
  /* fppowtf32.vhdl:1151:24  */
  assign n4464 = x == 10'b0000100001;
  /* fppowtf32.vhdl:1152:24  */
  assign n4467 = x == 10'b0000100010;
  /* fppowtf32.vhdl:1153:24  */
  assign n4470 = x == 10'b0000100011;
  /* fppowtf32.vhdl:1154:24  */
  assign n4473 = x == 10'b0000100100;
  /* fppowtf32.vhdl:1155:24  */
  assign n4476 = x == 10'b0000100101;
  /* fppowtf32.vhdl:1156:24  */
  assign n4479 = x == 10'b0000100110;
  /* fppowtf32.vhdl:1157:24  */
  assign n4482 = x == 10'b0000100111;
  /* fppowtf32.vhdl:1158:24  */
  assign n4485 = x == 10'b0000101000;
  /* fppowtf32.vhdl:1159:24  */
  assign n4488 = x == 10'b0000101001;
  /* fppowtf32.vhdl:1160:24  */
  assign n4491 = x == 10'b0000101010;
  /* fppowtf32.vhdl:1161:24  */
  assign n4494 = x == 10'b0000101011;
  /* fppowtf32.vhdl:1162:24  */
  assign n4497 = x == 10'b0000101100;
  /* fppowtf32.vhdl:1163:24  */
  assign n4500 = x == 10'b0000101101;
  /* fppowtf32.vhdl:1164:24  */
  assign n4503 = x == 10'b0000101110;
  /* fppowtf32.vhdl:1165:24  */
  assign n4506 = x == 10'b0000101111;
  /* fppowtf32.vhdl:1166:24  */
  assign n4509 = x == 10'b0000110000;
  /* fppowtf32.vhdl:1167:24  */
  assign n4512 = x == 10'b0000110001;
  /* fppowtf32.vhdl:1168:24  */
  assign n4515 = x == 10'b0000110010;
  /* fppowtf32.vhdl:1169:24  */
  assign n4518 = x == 10'b0000110011;
  /* fppowtf32.vhdl:1170:24  */
  assign n4521 = x == 10'b0000110100;
  /* fppowtf32.vhdl:1171:24  */
  assign n4524 = x == 10'b0000110101;
  /* fppowtf32.vhdl:1172:24  */
  assign n4527 = x == 10'b0000110110;
  /* fppowtf32.vhdl:1173:24  */
  assign n4530 = x == 10'b0000110111;
  /* fppowtf32.vhdl:1174:24  */
  assign n4533 = x == 10'b0000111000;
  /* fppowtf32.vhdl:1175:24  */
  assign n4536 = x == 10'b0000111001;
  /* fppowtf32.vhdl:1176:24  */
  assign n4539 = x == 10'b0000111010;
  /* fppowtf32.vhdl:1177:24  */
  assign n4542 = x == 10'b0000111011;
  /* fppowtf32.vhdl:1178:24  */
  assign n4545 = x == 10'b0000111100;
  /* fppowtf32.vhdl:1179:24  */
  assign n4548 = x == 10'b0000111101;
  /* fppowtf32.vhdl:1180:24  */
  assign n4551 = x == 10'b0000111110;
  /* fppowtf32.vhdl:1181:24  */
  assign n4554 = x == 10'b0000111111;
  /* fppowtf32.vhdl:1182:24  */
  assign n4557 = x == 10'b0001000000;
  /* fppowtf32.vhdl:1183:24  */
  assign n4560 = x == 10'b0001000001;
  /* fppowtf32.vhdl:1184:24  */
  assign n4563 = x == 10'b0001000010;
  /* fppowtf32.vhdl:1185:24  */
  assign n4566 = x == 10'b0001000011;
  /* fppowtf32.vhdl:1186:24  */
  assign n4569 = x == 10'b0001000100;
  /* fppowtf32.vhdl:1187:24  */
  assign n4572 = x == 10'b0001000101;
  /* fppowtf32.vhdl:1188:24  */
  assign n4575 = x == 10'b0001000110;
  /* fppowtf32.vhdl:1189:24  */
  assign n4578 = x == 10'b0001000111;
  /* fppowtf32.vhdl:1190:24  */
  assign n4581 = x == 10'b0001001000;
  /* fppowtf32.vhdl:1191:24  */
  assign n4584 = x == 10'b0001001001;
  /* fppowtf32.vhdl:1192:24  */
  assign n4587 = x == 10'b0001001010;
  /* fppowtf32.vhdl:1193:24  */
  assign n4590 = x == 10'b0001001011;
  /* fppowtf32.vhdl:1194:24  */
  assign n4593 = x == 10'b0001001100;
  /* fppowtf32.vhdl:1195:24  */
  assign n4596 = x == 10'b0001001101;
  /* fppowtf32.vhdl:1196:24  */
  assign n4599 = x == 10'b0001001110;
  /* fppowtf32.vhdl:1197:24  */
  assign n4602 = x == 10'b0001001111;
  /* fppowtf32.vhdl:1198:24  */
  assign n4605 = x == 10'b0001010000;
  /* fppowtf32.vhdl:1199:24  */
  assign n4608 = x == 10'b0001010001;
  /* fppowtf32.vhdl:1200:24  */
  assign n4611 = x == 10'b0001010010;
  /* fppowtf32.vhdl:1201:24  */
  assign n4614 = x == 10'b0001010011;
  /* fppowtf32.vhdl:1202:24  */
  assign n4617 = x == 10'b0001010100;
  /* fppowtf32.vhdl:1203:24  */
  assign n4620 = x == 10'b0001010101;
  /* fppowtf32.vhdl:1204:24  */
  assign n4623 = x == 10'b0001010110;
  /* fppowtf32.vhdl:1205:24  */
  assign n4626 = x == 10'b0001010111;
  /* fppowtf32.vhdl:1206:24  */
  assign n4629 = x == 10'b0001011000;
  /* fppowtf32.vhdl:1207:24  */
  assign n4632 = x == 10'b0001011001;
  /* fppowtf32.vhdl:1208:24  */
  assign n4635 = x == 10'b0001011010;
  /* fppowtf32.vhdl:1209:24  */
  assign n4638 = x == 10'b0001011011;
  /* fppowtf32.vhdl:1210:24  */
  assign n4641 = x == 10'b0001011100;
  /* fppowtf32.vhdl:1211:24  */
  assign n4644 = x == 10'b0001011101;
  /* fppowtf32.vhdl:1212:24  */
  assign n4647 = x == 10'b0001011110;
  /* fppowtf32.vhdl:1213:24  */
  assign n4650 = x == 10'b0001011111;
  /* fppowtf32.vhdl:1214:24  */
  assign n4653 = x == 10'b0001100000;
  /* fppowtf32.vhdl:1215:24  */
  assign n4656 = x == 10'b0001100001;
  /* fppowtf32.vhdl:1216:24  */
  assign n4659 = x == 10'b0001100010;
  /* fppowtf32.vhdl:1217:24  */
  assign n4662 = x == 10'b0001100011;
  /* fppowtf32.vhdl:1218:24  */
  assign n4665 = x == 10'b0001100100;
  /* fppowtf32.vhdl:1219:24  */
  assign n4668 = x == 10'b0001100101;
  /* fppowtf32.vhdl:1220:24  */
  assign n4671 = x == 10'b0001100110;
  /* fppowtf32.vhdl:1221:24  */
  assign n4674 = x == 10'b0001100111;
  /* fppowtf32.vhdl:1222:24  */
  assign n4677 = x == 10'b0001101000;
  /* fppowtf32.vhdl:1223:24  */
  assign n4680 = x == 10'b0001101001;
  /* fppowtf32.vhdl:1224:24  */
  assign n4683 = x == 10'b0001101010;
  /* fppowtf32.vhdl:1225:24  */
  assign n4686 = x == 10'b0001101011;
  /* fppowtf32.vhdl:1226:24  */
  assign n4689 = x == 10'b0001101100;
  /* fppowtf32.vhdl:1227:24  */
  assign n4692 = x == 10'b0001101101;
  /* fppowtf32.vhdl:1228:24  */
  assign n4695 = x == 10'b0001101110;
  /* fppowtf32.vhdl:1229:24  */
  assign n4698 = x == 10'b0001101111;
  /* fppowtf32.vhdl:1230:24  */
  assign n4701 = x == 10'b0001110000;
  /* fppowtf32.vhdl:1231:24  */
  assign n4704 = x == 10'b0001110001;
  /* fppowtf32.vhdl:1232:24  */
  assign n4707 = x == 10'b0001110010;
  /* fppowtf32.vhdl:1233:24  */
  assign n4710 = x == 10'b0001110011;
  /* fppowtf32.vhdl:1234:24  */
  assign n4713 = x == 10'b0001110100;
  /* fppowtf32.vhdl:1235:24  */
  assign n4716 = x == 10'b0001110101;
  /* fppowtf32.vhdl:1236:24  */
  assign n4719 = x == 10'b0001110110;
  /* fppowtf32.vhdl:1237:24  */
  assign n4722 = x == 10'b0001110111;
  /* fppowtf32.vhdl:1238:24  */
  assign n4725 = x == 10'b0001111000;
  /* fppowtf32.vhdl:1239:24  */
  assign n4728 = x == 10'b0001111001;
  /* fppowtf32.vhdl:1240:24  */
  assign n4731 = x == 10'b0001111010;
  /* fppowtf32.vhdl:1241:24  */
  assign n4734 = x == 10'b0001111011;
  /* fppowtf32.vhdl:1242:24  */
  assign n4737 = x == 10'b0001111100;
  /* fppowtf32.vhdl:1243:24  */
  assign n4740 = x == 10'b0001111101;
  /* fppowtf32.vhdl:1244:24  */
  assign n4743 = x == 10'b0001111110;
  /* fppowtf32.vhdl:1245:24  */
  assign n4746 = x == 10'b0001111111;
  /* fppowtf32.vhdl:1246:24  */
  assign n4749 = x == 10'b0010000000;
  /* fppowtf32.vhdl:1247:24  */
  assign n4752 = x == 10'b0010000001;
  /* fppowtf32.vhdl:1248:24  */
  assign n4755 = x == 10'b0010000010;
  /* fppowtf32.vhdl:1249:24  */
  assign n4758 = x == 10'b0010000011;
  /* fppowtf32.vhdl:1250:24  */
  assign n4761 = x == 10'b0010000100;
  /* fppowtf32.vhdl:1251:24  */
  assign n4764 = x == 10'b0010000101;
  /* fppowtf32.vhdl:1252:24  */
  assign n4767 = x == 10'b0010000110;
  /* fppowtf32.vhdl:1253:24  */
  assign n4770 = x == 10'b0010000111;
  /* fppowtf32.vhdl:1254:24  */
  assign n4773 = x == 10'b0010001000;
  /* fppowtf32.vhdl:1255:24  */
  assign n4776 = x == 10'b0010001001;
  /* fppowtf32.vhdl:1256:24  */
  assign n4779 = x == 10'b0010001010;
  /* fppowtf32.vhdl:1257:24  */
  assign n4782 = x == 10'b0010001011;
  /* fppowtf32.vhdl:1258:24  */
  assign n4785 = x == 10'b0010001100;
  /* fppowtf32.vhdl:1259:24  */
  assign n4788 = x == 10'b0010001101;
  /* fppowtf32.vhdl:1260:24  */
  assign n4791 = x == 10'b0010001110;
  /* fppowtf32.vhdl:1261:24  */
  assign n4794 = x == 10'b0010001111;
  /* fppowtf32.vhdl:1262:24  */
  assign n4797 = x == 10'b0010010000;
  /* fppowtf32.vhdl:1263:24  */
  assign n4800 = x == 10'b0010010001;
  /* fppowtf32.vhdl:1264:24  */
  assign n4803 = x == 10'b0010010010;
  /* fppowtf32.vhdl:1265:24  */
  assign n4806 = x == 10'b0010010011;
  /* fppowtf32.vhdl:1266:24  */
  assign n4809 = x == 10'b0010010100;
  /* fppowtf32.vhdl:1267:24  */
  assign n4812 = x == 10'b0010010101;
  /* fppowtf32.vhdl:1268:24  */
  assign n4815 = x == 10'b0010010110;
  /* fppowtf32.vhdl:1269:24  */
  assign n4818 = x == 10'b0010010111;
  /* fppowtf32.vhdl:1270:24  */
  assign n4821 = x == 10'b0010011000;
  /* fppowtf32.vhdl:1271:24  */
  assign n4824 = x == 10'b0010011001;
  /* fppowtf32.vhdl:1272:24  */
  assign n4827 = x == 10'b0010011010;
  /* fppowtf32.vhdl:1273:24  */
  assign n4830 = x == 10'b0010011011;
  /* fppowtf32.vhdl:1274:24  */
  assign n4833 = x == 10'b0010011100;
  /* fppowtf32.vhdl:1275:24  */
  assign n4836 = x == 10'b0010011101;
  /* fppowtf32.vhdl:1276:24  */
  assign n4839 = x == 10'b0010011110;
  /* fppowtf32.vhdl:1277:24  */
  assign n4842 = x == 10'b0010011111;
  /* fppowtf32.vhdl:1278:24  */
  assign n4845 = x == 10'b0010100000;
  /* fppowtf32.vhdl:1279:24  */
  assign n4848 = x == 10'b0010100001;
  /* fppowtf32.vhdl:1280:24  */
  assign n4851 = x == 10'b0010100010;
  /* fppowtf32.vhdl:1281:24  */
  assign n4854 = x == 10'b0010100011;
  /* fppowtf32.vhdl:1282:24  */
  assign n4857 = x == 10'b0010100100;
  /* fppowtf32.vhdl:1283:24  */
  assign n4860 = x == 10'b0010100101;
  /* fppowtf32.vhdl:1284:24  */
  assign n4863 = x == 10'b0010100110;
  /* fppowtf32.vhdl:1285:24  */
  assign n4866 = x == 10'b0010100111;
  /* fppowtf32.vhdl:1286:24  */
  assign n4869 = x == 10'b0010101000;
  /* fppowtf32.vhdl:1287:24  */
  assign n4872 = x == 10'b0010101001;
  /* fppowtf32.vhdl:1288:24  */
  assign n4875 = x == 10'b0010101010;
  /* fppowtf32.vhdl:1289:24  */
  assign n4878 = x == 10'b0010101011;
  /* fppowtf32.vhdl:1290:24  */
  assign n4881 = x == 10'b0010101100;
  /* fppowtf32.vhdl:1291:24  */
  assign n4884 = x == 10'b0010101101;
  /* fppowtf32.vhdl:1292:24  */
  assign n4887 = x == 10'b0010101110;
  /* fppowtf32.vhdl:1293:24  */
  assign n4890 = x == 10'b0010101111;
  /* fppowtf32.vhdl:1294:24  */
  assign n4893 = x == 10'b0010110000;
  /* fppowtf32.vhdl:1295:24  */
  assign n4896 = x == 10'b0010110001;
  /* fppowtf32.vhdl:1296:24  */
  assign n4899 = x == 10'b0010110010;
  /* fppowtf32.vhdl:1297:24  */
  assign n4902 = x == 10'b0010110011;
  /* fppowtf32.vhdl:1298:24  */
  assign n4905 = x == 10'b0010110100;
  /* fppowtf32.vhdl:1299:24  */
  assign n4908 = x == 10'b0010110101;
  /* fppowtf32.vhdl:1300:24  */
  assign n4911 = x == 10'b0010110110;
  /* fppowtf32.vhdl:1301:24  */
  assign n4914 = x == 10'b0010110111;
  /* fppowtf32.vhdl:1302:24  */
  assign n4917 = x == 10'b0010111000;
  /* fppowtf32.vhdl:1303:24  */
  assign n4920 = x == 10'b0010111001;
  /* fppowtf32.vhdl:1304:24  */
  assign n4923 = x == 10'b0010111010;
  /* fppowtf32.vhdl:1305:24  */
  assign n4926 = x == 10'b0010111011;
  /* fppowtf32.vhdl:1306:24  */
  assign n4929 = x == 10'b0010111100;
  /* fppowtf32.vhdl:1307:24  */
  assign n4932 = x == 10'b0010111101;
  /* fppowtf32.vhdl:1308:24  */
  assign n4935 = x == 10'b0010111110;
  /* fppowtf32.vhdl:1309:24  */
  assign n4938 = x == 10'b0010111111;
  /* fppowtf32.vhdl:1310:24  */
  assign n4941 = x == 10'b0011000000;
  /* fppowtf32.vhdl:1311:24  */
  assign n4944 = x == 10'b0011000001;
  /* fppowtf32.vhdl:1312:24  */
  assign n4947 = x == 10'b0011000010;
  /* fppowtf32.vhdl:1313:24  */
  assign n4950 = x == 10'b0011000011;
  /* fppowtf32.vhdl:1314:24  */
  assign n4953 = x == 10'b0011000100;
  /* fppowtf32.vhdl:1315:24  */
  assign n4956 = x == 10'b0011000101;
  /* fppowtf32.vhdl:1316:24  */
  assign n4959 = x == 10'b0011000110;
  /* fppowtf32.vhdl:1317:24  */
  assign n4962 = x == 10'b0011000111;
  /* fppowtf32.vhdl:1318:24  */
  assign n4965 = x == 10'b0011001000;
  /* fppowtf32.vhdl:1319:24  */
  assign n4968 = x == 10'b0011001001;
  /* fppowtf32.vhdl:1320:24  */
  assign n4971 = x == 10'b0011001010;
  /* fppowtf32.vhdl:1321:24  */
  assign n4974 = x == 10'b0011001011;
  /* fppowtf32.vhdl:1322:24  */
  assign n4977 = x == 10'b0011001100;
  /* fppowtf32.vhdl:1323:24  */
  assign n4980 = x == 10'b0011001101;
  /* fppowtf32.vhdl:1324:24  */
  assign n4983 = x == 10'b0011001110;
  /* fppowtf32.vhdl:1325:24  */
  assign n4986 = x == 10'b0011001111;
  /* fppowtf32.vhdl:1326:24  */
  assign n4989 = x == 10'b0011010000;
  /* fppowtf32.vhdl:1327:24  */
  assign n4992 = x == 10'b0011010001;
  /* fppowtf32.vhdl:1328:24  */
  assign n4995 = x == 10'b0011010010;
  /* fppowtf32.vhdl:1329:24  */
  assign n4998 = x == 10'b0011010011;
  /* fppowtf32.vhdl:1330:24  */
  assign n5001 = x == 10'b0011010100;
  /* fppowtf32.vhdl:1331:24  */
  assign n5004 = x == 10'b0011010101;
  /* fppowtf32.vhdl:1332:24  */
  assign n5007 = x == 10'b0011010110;
  /* fppowtf32.vhdl:1333:24  */
  assign n5010 = x == 10'b0011010111;
  /* fppowtf32.vhdl:1334:24  */
  assign n5013 = x == 10'b0011011000;
  /* fppowtf32.vhdl:1335:24  */
  assign n5016 = x == 10'b0011011001;
  /* fppowtf32.vhdl:1336:24  */
  assign n5019 = x == 10'b0011011010;
  /* fppowtf32.vhdl:1337:24  */
  assign n5022 = x == 10'b0011011011;
  /* fppowtf32.vhdl:1338:24  */
  assign n5025 = x == 10'b0011011100;
  /* fppowtf32.vhdl:1339:24  */
  assign n5028 = x == 10'b0011011101;
  /* fppowtf32.vhdl:1340:24  */
  assign n5031 = x == 10'b0011011110;
  /* fppowtf32.vhdl:1341:24  */
  assign n5034 = x == 10'b0011011111;
  /* fppowtf32.vhdl:1342:24  */
  assign n5037 = x == 10'b0011100000;
  /* fppowtf32.vhdl:1343:24  */
  assign n5040 = x == 10'b0011100001;
  /* fppowtf32.vhdl:1344:24  */
  assign n5043 = x == 10'b0011100010;
  /* fppowtf32.vhdl:1345:24  */
  assign n5046 = x == 10'b0011100011;
  /* fppowtf32.vhdl:1346:24  */
  assign n5049 = x == 10'b0011100100;
  /* fppowtf32.vhdl:1347:24  */
  assign n5052 = x == 10'b0011100101;
  /* fppowtf32.vhdl:1348:24  */
  assign n5055 = x == 10'b0011100110;
  /* fppowtf32.vhdl:1349:24  */
  assign n5058 = x == 10'b0011100111;
  /* fppowtf32.vhdl:1350:24  */
  assign n5061 = x == 10'b0011101000;
  /* fppowtf32.vhdl:1351:24  */
  assign n5064 = x == 10'b0011101001;
  /* fppowtf32.vhdl:1352:24  */
  assign n5067 = x == 10'b0011101010;
  /* fppowtf32.vhdl:1353:24  */
  assign n5070 = x == 10'b0011101011;
  /* fppowtf32.vhdl:1354:24  */
  assign n5073 = x == 10'b0011101100;
  /* fppowtf32.vhdl:1355:24  */
  assign n5076 = x == 10'b0011101101;
  /* fppowtf32.vhdl:1356:24  */
  assign n5079 = x == 10'b0011101110;
  /* fppowtf32.vhdl:1357:24  */
  assign n5082 = x == 10'b0011101111;
  /* fppowtf32.vhdl:1358:24  */
  assign n5085 = x == 10'b0011110000;
  /* fppowtf32.vhdl:1359:24  */
  assign n5088 = x == 10'b0011110001;
  /* fppowtf32.vhdl:1360:24  */
  assign n5091 = x == 10'b0011110010;
  /* fppowtf32.vhdl:1361:24  */
  assign n5094 = x == 10'b0011110011;
  /* fppowtf32.vhdl:1362:24  */
  assign n5097 = x == 10'b0011110100;
  /* fppowtf32.vhdl:1363:24  */
  assign n5100 = x == 10'b0011110101;
  /* fppowtf32.vhdl:1364:24  */
  assign n5103 = x == 10'b0011110110;
  /* fppowtf32.vhdl:1365:24  */
  assign n5106 = x == 10'b0011110111;
  /* fppowtf32.vhdl:1366:24  */
  assign n5109 = x == 10'b0011111000;
  /* fppowtf32.vhdl:1367:24  */
  assign n5112 = x == 10'b0011111001;
  /* fppowtf32.vhdl:1368:24  */
  assign n5115 = x == 10'b0011111010;
  /* fppowtf32.vhdl:1369:24  */
  assign n5118 = x == 10'b0011111011;
  /* fppowtf32.vhdl:1370:24  */
  assign n5121 = x == 10'b0011111100;
  /* fppowtf32.vhdl:1371:24  */
  assign n5124 = x == 10'b0011111101;
  /* fppowtf32.vhdl:1372:24  */
  assign n5127 = x == 10'b0011111110;
  /* fppowtf32.vhdl:1373:24  */
  assign n5130 = x == 10'b0011111111;
  /* fppowtf32.vhdl:1374:24  */
  assign n5133 = x == 10'b0100000000;
  /* fppowtf32.vhdl:1375:24  */
  assign n5136 = x == 10'b0100000001;
  /* fppowtf32.vhdl:1376:24  */
  assign n5139 = x == 10'b0100000010;
  /* fppowtf32.vhdl:1377:24  */
  assign n5142 = x == 10'b0100000011;
  /* fppowtf32.vhdl:1378:24  */
  assign n5145 = x == 10'b0100000100;
  /* fppowtf32.vhdl:1379:24  */
  assign n5148 = x == 10'b0100000101;
  /* fppowtf32.vhdl:1380:24  */
  assign n5151 = x == 10'b0100000110;
  /* fppowtf32.vhdl:1381:24  */
  assign n5154 = x == 10'b0100000111;
  /* fppowtf32.vhdl:1382:24  */
  assign n5157 = x == 10'b0100001000;
  /* fppowtf32.vhdl:1383:24  */
  assign n5160 = x == 10'b0100001001;
  /* fppowtf32.vhdl:1384:24  */
  assign n5163 = x == 10'b0100001010;
  /* fppowtf32.vhdl:1385:24  */
  assign n5166 = x == 10'b0100001011;
  /* fppowtf32.vhdl:1386:24  */
  assign n5169 = x == 10'b0100001100;
  /* fppowtf32.vhdl:1387:24  */
  assign n5172 = x == 10'b0100001101;
  /* fppowtf32.vhdl:1388:24  */
  assign n5175 = x == 10'b0100001110;
  /* fppowtf32.vhdl:1389:24  */
  assign n5178 = x == 10'b0100001111;
  /* fppowtf32.vhdl:1390:24  */
  assign n5181 = x == 10'b0100010000;
  /* fppowtf32.vhdl:1391:24  */
  assign n5184 = x == 10'b0100010001;
  /* fppowtf32.vhdl:1392:24  */
  assign n5187 = x == 10'b0100010010;
  /* fppowtf32.vhdl:1393:24  */
  assign n5190 = x == 10'b0100010011;
  /* fppowtf32.vhdl:1394:24  */
  assign n5193 = x == 10'b0100010100;
  /* fppowtf32.vhdl:1395:24  */
  assign n5196 = x == 10'b0100010101;
  /* fppowtf32.vhdl:1396:24  */
  assign n5199 = x == 10'b0100010110;
  /* fppowtf32.vhdl:1397:24  */
  assign n5202 = x == 10'b0100010111;
  /* fppowtf32.vhdl:1398:24  */
  assign n5205 = x == 10'b0100011000;
  /* fppowtf32.vhdl:1399:24  */
  assign n5208 = x == 10'b0100011001;
  /* fppowtf32.vhdl:1400:24  */
  assign n5211 = x == 10'b0100011010;
  /* fppowtf32.vhdl:1401:24  */
  assign n5214 = x == 10'b0100011011;
  /* fppowtf32.vhdl:1402:24  */
  assign n5217 = x == 10'b0100011100;
  /* fppowtf32.vhdl:1403:24  */
  assign n5220 = x == 10'b0100011101;
  /* fppowtf32.vhdl:1404:24  */
  assign n5223 = x == 10'b0100011110;
  /* fppowtf32.vhdl:1405:24  */
  assign n5226 = x == 10'b0100011111;
  /* fppowtf32.vhdl:1406:24  */
  assign n5229 = x == 10'b0100100000;
  /* fppowtf32.vhdl:1407:24  */
  assign n5232 = x == 10'b0100100001;
  /* fppowtf32.vhdl:1408:24  */
  assign n5235 = x == 10'b0100100010;
  /* fppowtf32.vhdl:1409:24  */
  assign n5238 = x == 10'b0100100011;
  /* fppowtf32.vhdl:1410:24  */
  assign n5241 = x == 10'b0100100100;
  /* fppowtf32.vhdl:1411:24  */
  assign n5244 = x == 10'b0100100101;
  /* fppowtf32.vhdl:1412:24  */
  assign n5247 = x == 10'b0100100110;
  /* fppowtf32.vhdl:1413:24  */
  assign n5250 = x == 10'b0100100111;
  /* fppowtf32.vhdl:1414:24  */
  assign n5253 = x == 10'b0100101000;
  /* fppowtf32.vhdl:1415:24  */
  assign n5256 = x == 10'b0100101001;
  /* fppowtf32.vhdl:1416:24  */
  assign n5259 = x == 10'b0100101010;
  /* fppowtf32.vhdl:1417:24  */
  assign n5262 = x == 10'b0100101011;
  /* fppowtf32.vhdl:1418:24  */
  assign n5265 = x == 10'b0100101100;
  /* fppowtf32.vhdl:1419:24  */
  assign n5268 = x == 10'b0100101101;
  /* fppowtf32.vhdl:1420:24  */
  assign n5271 = x == 10'b0100101110;
  /* fppowtf32.vhdl:1421:24  */
  assign n5274 = x == 10'b0100101111;
  /* fppowtf32.vhdl:1422:24  */
  assign n5277 = x == 10'b0100110000;
  /* fppowtf32.vhdl:1423:24  */
  assign n5280 = x == 10'b0100110001;
  /* fppowtf32.vhdl:1424:24  */
  assign n5283 = x == 10'b0100110010;
  /* fppowtf32.vhdl:1425:24  */
  assign n5286 = x == 10'b0100110011;
  /* fppowtf32.vhdl:1426:24  */
  assign n5289 = x == 10'b0100110100;
  /* fppowtf32.vhdl:1427:24  */
  assign n5292 = x == 10'b0100110101;
  /* fppowtf32.vhdl:1428:24  */
  assign n5295 = x == 10'b0100110110;
  /* fppowtf32.vhdl:1429:24  */
  assign n5298 = x == 10'b0100110111;
  /* fppowtf32.vhdl:1430:24  */
  assign n5301 = x == 10'b0100111000;
  /* fppowtf32.vhdl:1431:24  */
  assign n5304 = x == 10'b0100111001;
  /* fppowtf32.vhdl:1432:24  */
  assign n5307 = x == 10'b0100111010;
  /* fppowtf32.vhdl:1433:24  */
  assign n5310 = x == 10'b0100111011;
  /* fppowtf32.vhdl:1434:24  */
  assign n5313 = x == 10'b0100111100;
  /* fppowtf32.vhdl:1435:24  */
  assign n5316 = x == 10'b0100111101;
  /* fppowtf32.vhdl:1436:24  */
  assign n5319 = x == 10'b0100111110;
  /* fppowtf32.vhdl:1437:24  */
  assign n5322 = x == 10'b0100111111;
  /* fppowtf32.vhdl:1438:24  */
  assign n5325 = x == 10'b0101000000;
  /* fppowtf32.vhdl:1439:24  */
  assign n5328 = x == 10'b0101000001;
  /* fppowtf32.vhdl:1440:24  */
  assign n5331 = x == 10'b0101000010;
  /* fppowtf32.vhdl:1441:24  */
  assign n5334 = x == 10'b0101000011;
  /* fppowtf32.vhdl:1442:24  */
  assign n5337 = x == 10'b0101000100;
  /* fppowtf32.vhdl:1443:24  */
  assign n5340 = x == 10'b0101000101;
  /* fppowtf32.vhdl:1444:24  */
  assign n5343 = x == 10'b0101000110;
  /* fppowtf32.vhdl:1445:24  */
  assign n5346 = x == 10'b0101000111;
  /* fppowtf32.vhdl:1446:24  */
  assign n5349 = x == 10'b0101001000;
  /* fppowtf32.vhdl:1447:24  */
  assign n5352 = x == 10'b0101001001;
  /* fppowtf32.vhdl:1448:24  */
  assign n5355 = x == 10'b0101001010;
  /* fppowtf32.vhdl:1449:24  */
  assign n5358 = x == 10'b0101001011;
  /* fppowtf32.vhdl:1450:24  */
  assign n5361 = x == 10'b0101001100;
  /* fppowtf32.vhdl:1451:24  */
  assign n5364 = x == 10'b0101001101;
  /* fppowtf32.vhdl:1452:24  */
  assign n5367 = x == 10'b0101001110;
  /* fppowtf32.vhdl:1453:24  */
  assign n5370 = x == 10'b0101001111;
  /* fppowtf32.vhdl:1454:24  */
  assign n5373 = x == 10'b0101010000;
  /* fppowtf32.vhdl:1455:24  */
  assign n5376 = x == 10'b0101010001;
  /* fppowtf32.vhdl:1456:24  */
  assign n5379 = x == 10'b0101010010;
  /* fppowtf32.vhdl:1457:24  */
  assign n5382 = x == 10'b0101010011;
  /* fppowtf32.vhdl:1458:24  */
  assign n5385 = x == 10'b0101010100;
  /* fppowtf32.vhdl:1459:24  */
  assign n5388 = x == 10'b0101010101;
  /* fppowtf32.vhdl:1460:24  */
  assign n5391 = x == 10'b0101010110;
  /* fppowtf32.vhdl:1461:24  */
  assign n5394 = x == 10'b0101010111;
  /* fppowtf32.vhdl:1462:24  */
  assign n5397 = x == 10'b0101011000;
  /* fppowtf32.vhdl:1463:24  */
  assign n5400 = x == 10'b0101011001;
  /* fppowtf32.vhdl:1464:24  */
  assign n5403 = x == 10'b0101011010;
  /* fppowtf32.vhdl:1465:24  */
  assign n5406 = x == 10'b0101011011;
  /* fppowtf32.vhdl:1466:24  */
  assign n5409 = x == 10'b0101011100;
  /* fppowtf32.vhdl:1467:24  */
  assign n5412 = x == 10'b0101011101;
  /* fppowtf32.vhdl:1468:24  */
  assign n5415 = x == 10'b0101011110;
  /* fppowtf32.vhdl:1469:24  */
  assign n5418 = x == 10'b0101011111;
  /* fppowtf32.vhdl:1470:24  */
  assign n5421 = x == 10'b0101100000;
  /* fppowtf32.vhdl:1471:24  */
  assign n5424 = x == 10'b0101100001;
  /* fppowtf32.vhdl:1472:24  */
  assign n5427 = x == 10'b0101100010;
  /* fppowtf32.vhdl:1473:24  */
  assign n5430 = x == 10'b0101100011;
  /* fppowtf32.vhdl:1474:24  */
  assign n5433 = x == 10'b0101100100;
  /* fppowtf32.vhdl:1475:24  */
  assign n5436 = x == 10'b0101100101;
  /* fppowtf32.vhdl:1476:24  */
  assign n5439 = x == 10'b0101100110;
  /* fppowtf32.vhdl:1477:24  */
  assign n5442 = x == 10'b0101100111;
  /* fppowtf32.vhdl:1478:24  */
  assign n5445 = x == 10'b0101101000;
  /* fppowtf32.vhdl:1479:24  */
  assign n5448 = x == 10'b0101101001;
  /* fppowtf32.vhdl:1480:24  */
  assign n5451 = x == 10'b0101101010;
  /* fppowtf32.vhdl:1481:24  */
  assign n5454 = x == 10'b0101101011;
  /* fppowtf32.vhdl:1482:24  */
  assign n5457 = x == 10'b0101101100;
  /* fppowtf32.vhdl:1483:24  */
  assign n5460 = x == 10'b0101101101;
  /* fppowtf32.vhdl:1484:24  */
  assign n5463 = x == 10'b0101101110;
  /* fppowtf32.vhdl:1485:24  */
  assign n5466 = x == 10'b0101101111;
  /* fppowtf32.vhdl:1486:24  */
  assign n5469 = x == 10'b0101110000;
  /* fppowtf32.vhdl:1487:24  */
  assign n5472 = x == 10'b0101110001;
  /* fppowtf32.vhdl:1488:24  */
  assign n5475 = x == 10'b0101110010;
  /* fppowtf32.vhdl:1489:24  */
  assign n5478 = x == 10'b0101110011;
  /* fppowtf32.vhdl:1490:24  */
  assign n5481 = x == 10'b0101110100;
  /* fppowtf32.vhdl:1491:24  */
  assign n5484 = x == 10'b0101110101;
  /* fppowtf32.vhdl:1492:24  */
  assign n5487 = x == 10'b0101110110;
  /* fppowtf32.vhdl:1493:24  */
  assign n5490 = x == 10'b0101110111;
  /* fppowtf32.vhdl:1494:24  */
  assign n5493 = x == 10'b0101111000;
  /* fppowtf32.vhdl:1495:24  */
  assign n5496 = x == 10'b0101111001;
  /* fppowtf32.vhdl:1496:24  */
  assign n5499 = x == 10'b0101111010;
  /* fppowtf32.vhdl:1497:24  */
  assign n5502 = x == 10'b0101111011;
  /* fppowtf32.vhdl:1498:24  */
  assign n5505 = x == 10'b0101111100;
  /* fppowtf32.vhdl:1499:24  */
  assign n5508 = x == 10'b0101111101;
  /* fppowtf32.vhdl:1500:24  */
  assign n5511 = x == 10'b0101111110;
  /* fppowtf32.vhdl:1501:24  */
  assign n5514 = x == 10'b0101111111;
  /* fppowtf32.vhdl:1502:24  */
  assign n5517 = x == 10'b0110000000;
  /* fppowtf32.vhdl:1503:24  */
  assign n5520 = x == 10'b0110000001;
  /* fppowtf32.vhdl:1504:24  */
  assign n5523 = x == 10'b0110000010;
  /* fppowtf32.vhdl:1505:24  */
  assign n5526 = x == 10'b0110000011;
  /* fppowtf32.vhdl:1506:24  */
  assign n5529 = x == 10'b0110000100;
  /* fppowtf32.vhdl:1507:24  */
  assign n5532 = x == 10'b0110000101;
  /* fppowtf32.vhdl:1508:24  */
  assign n5535 = x == 10'b0110000110;
  /* fppowtf32.vhdl:1509:24  */
  assign n5538 = x == 10'b0110000111;
  /* fppowtf32.vhdl:1510:24  */
  assign n5541 = x == 10'b0110001000;
  /* fppowtf32.vhdl:1511:24  */
  assign n5544 = x == 10'b0110001001;
  /* fppowtf32.vhdl:1512:24  */
  assign n5547 = x == 10'b0110001010;
  /* fppowtf32.vhdl:1513:24  */
  assign n5550 = x == 10'b0110001011;
  /* fppowtf32.vhdl:1514:24  */
  assign n5553 = x == 10'b0110001100;
  /* fppowtf32.vhdl:1515:24  */
  assign n5556 = x == 10'b0110001101;
  /* fppowtf32.vhdl:1516:24  */
  assign n5559 = x == 10'b0110001110;
  /* fppowtf32.vhdl:1517:24  */
  assign n5562 = x == 10'b0110001111;
  /* fppowtf32.vhdl:1518:24  */
  assign n5565 = x == 10'b0110010000;
  /* fppowtf32.vhdl:1519:24  */
  assign n5568 = x == 10'b0110010001;
  /* fppowtf32.vhdl:1520:24  */
  assign n5571 = x == 10'b0110010010;
  /* fppowtf32.vhdl:1521:24  */
  assign n5574 = x == 10'b0110010011;
  /* fppowtf32.vhdl:1522:24  */
  assign n5577 = x == 10'b0110010100;
  /* fppowtf32.vhdl:1523:24  */
  assign n5580 = x == 10'b0110010101;
  /* fppowtf32.vhdl:1524:24  */
  assign n5583 = x == 10'b0110010110;
  /* fppowtf32.vhdl:1525:24  */
  assign n5586 = x == 10'b0110010111;
  /* fppowtf32.vhdl:1526:24  */
  assign n5589 = x == 10'b0110011000;
  /* fppowtf32.vhdl:1527:24  */
  assign n5592 = x == 10'b0110011001;
  /* fppowtf32.vhdl:1528:24  */
  assign n5595 = x == 10'b0110011010;
  /* fppowtf32.vhdl:1529:24  */
  assign n5598 = x == 10'b0110011011;
  /* fppowtf32.vhdl:1530:24  */
  assign n5601 = x == 10'b0110011100;
  /* fppowtf32.vhdl:1531:24  */
  assign n5604 = x == 10'b0110011101;
  /* fppowtf32.vhdl:1532:24  */
  assign n5607 = x == 10'b0110011110;
  /* fppowtf32.vhdl:1533:24  */
  assign n5610 = x == 10'b0110011111;
  /* fppowtf32.vhdl:1534:24  */
  assign n5613 = x == 10'b0110100000;
  /* fppowtf32.vhdl:1535:24  */
  assign n5616 = x == 10'b0110100001;
  /* fppowtf32.vhdl:1536:24  */
  assign n5619 = x == 10'b0110100010;
  /* fppowtf32.vhdl:1537:24  */
  assign n5622 = x == 10'b0110100011;
  /* fppowtf32.vhdl:1538:24  */
  assign n5625 = x == 10'b0110100100;
  /* fppowtf32.vhdl:1539:24  */
  assign n5628 = x == 10'b0110100101;
  /* fppowtf32.vhdl:1540:24  */
  assign n5631 = x == 10'b0110100110;
  /* fppowtf32.vhdl:1541:24  */
  assign n5634 = x == 10'b0110100111;
  /* fppowtf32.vhdl:1542:24  */
  assign n5637 = x == 10'b0110101000;
  /* fppowtf32.vhdl:1543:24  */
  assign n5640 = x == 10'b0110101001;
  /* fppowtf32.vhdl:1544:24  */
  assign n5643 = x == 10'b0110101010;
  /* fppowtf32.vhdl:1545:24  */
  assign n5646 = x == 10'b0110101011;
  /* fppowtf32.vhdl:1546:24  */
  assign n5649 = x == 10'b0110101100;
  /* fppowtf32.vhdl:1547:24  */
  assign n5652 = x == 10'b0110101101;
  /* fppowtf32.vhdl:1548:24  */
  assign n5655 = x == 10'b0110101110;
  /* fppowtf32.vhdl:1549:24  */
  assign n5658 = x == 10'b0110101111;
  /* fppowtf32.vhdl:1550:24  */
  assign n5661 = x == 10'b0110110000;
  /* fppowtf32.vhdl:1551:24  */
  assign n5664 = x == 10'b0110110001;
  /* fppowtf32.vhdl:1552:24  */
  assign n5667 = x == 10'b0110110010;
  /* fppowtf32.vhdl:1553:24  */
  assign n5670 = x == 10'b0110110011;
  /* fppowtf32.vhdl:1554:24  */
  assign n5673 = x == 10'b0110110100;
  /* fppowtf32.vhdl:1555:24  */
  assign n5676 = x == 10'b0110110101;
  /* fppowtf32.vhdl:1556:24  */
  assign n5679 = x == 10'b0110110110;
  /* fppowtf32.vhdl:1557:24  */
  assign n5682 = x == 10'b0110110111;
  /* fppowtf32.vhdl:1558:24  */
  assign n5685 = x == 10'b0110111000;
  /* fppowtf32.vhdl:1559:24  */
  assign n5688 = x == 10'b0110111001;
  /* fppowtf32.vhdl:1560:24  */
  assign n5691 = x == 10'b0110111010;
  /* fppowtf32.vhdl:1561:24  */
  assign n5694 = x == 10'b0110111011;
  /* fppowtf32.vhdl:1562:24  */
  assign n5697 = x == 10'b0110111100;
  /* fppowtf32.vhdl:1563:24  */
  assign n5700 = x == 10'b0110111101;
  /* fppowtf32.vhdl:1564:24  */
  assign n5703 = x == 10'b0110111110;
  /* fppowtf32.vhdl:1565:24  */
  assign n5706 = x == 10'b0110111111;
  /* fppowtf32.vhdl:1566:24  */
  assign n5709 = x == 10'b0111000000;
  /* fppowtf32.vhdl:1567:24  */
  assign n5712 = x == 10'b0111000001;
  /* fppowtf32.vhdl:1568:24  */
  assign n5715 = x == 10'b0111000010;
  /* fppowtf32.vhdl:1569:24  */
  assign n5718 = x == 10'b0111000011;
  /* fppowtf32.vhdl:1570:24  */
  assign n5721 = x == 10'b0111000100;
  /* fppowtf32.vhdl:1571:24  */
  assign n5724 = x == 10'b0111000101;
  /* fppowtf32.vhdl:1572:24  */
  assign n5727 = x == 10'b0111000110;
  /* fppowtf32.vhdl:1573:24  */
  assign n5730 = x == 10'b0111000111;
  /* fppowtf32.vhdl:1574:24  */
  assign n5733 = x == 10'b0111001000;
  /* fppowtf32.vhdl:1575:24  */
  assign n5736 = x == 10'b0111001001;
  /* fppowtf32.vhdl:1576:24  */
  assign n5739 = x == 10'b0111001010;
  /* fppowtf32.vhdl:1577:24  */
  assign n5742 = x == 10'b0111001011;
  /* fppowtf32.vhdl:1578:24  */
  assign n5745 = x == 10'b0111001100;
  /* fppowtf32.vhdl:1579:24  */
  assign n5748 = x == 10'b0111001101;
  /* fppowtf32.vhdl:1580:24  */
  assign n5751 = x == 10'b0111001110;
  /* fppowtf32.vhdl:1581:24  */
  assign n5754 = x == 10'b0111001111;
  /* fppowtf32.vhdl:1582:24  */
  assign n5757 = x == 10'b0111010000;
  /* fppowtf32.vhdl:1583:24  */
  assign n5760 = x == 10'b0111010001;
  /* fppowtf32.vhdl:1584:24  */
  assign n5763 = x == 10'b0111010010;
  /* fppowtf32.vhdl:1585:24  */
  assign n5766 = x == 10'b0111010011;
  /* fppowtf32.vhdl:1586:24  */
  assign n5769 = x == 10'b0111010100;
  /* fppowtf32.vhdl:1587:24  */
  assign n5772 = x == 10'b0111010101;
  /* fppowtf32.vhdl:1588:24  */
  assign n5775 = x == 10'b0111010110;
  /* fppowtf32.vhdl:1589:24  */
  assign n5778 = x == 10'b0111010111;
  /* fppowtf32.vhdl:1590:24  */
  assign n5781 = x == 10'b0111011000;
  /* fppowtf32.vhdl:1591:24  */
  assign n5784 = x == 10'b0111011001;
  /* fppowtf32.vhdl:1592:24  */
  assign n5787 = x == 10'b0111011010;
  /* fppowtf32.vhdl:1593:24  */
  assign n5790 = x == 10'b0111011011;
  /* fppowtf32.vhdl:1594:24  */
  assign n5793 = x == 10'b0111011100;
  /* fppowtf32.vhdl:1595:24  */
  assign n5796 = x == 10'b0111011101;
  /* fppowtf32.vhdl:1596:24  */
  assign n5799 = x == 10'b0111011110;
  /* fppowtf32.vhdl:1597:24  */
  assign n5802 = x == 10'b0111011111;
  /* fppowtf32.vhdl:1598:24  */
  assign n5805 = x == 10'b0111100000;
  /* fppowtf32.vhdl:1599:24  */
  assign n5808 = x == 10'b0111100001;
  /* fppowtf32.vhdl:1600:24  */
  assign n5811 = x == 10'b0111100010;
  /* fppowtf32.vhdl:1601:24  */
  assign n5814 = x == 10'b0111100011;
  /* fppowtf32.vhdl:1602:24  */
  assign n5817 = x == 10'b0111100100;
  /* fppowtf32.vhdl:1603:24  */
  assign n5820 = x == 10'b0111100101;
  /* fppowtf32.vhdl:1604:24  */
  assign n5823 = x == 10'b0111100110;
  /* fppowtf32.vhdl:1605:24  */
  assign n5826 = x == 10'b0111100111;
  /* fppowtf32.vhdl:1606:24  */
  assign n5829 = x == 10'b0111101000;
  /* fppowtf32.vhdl:1607:24  */
  assign n5832 = x == 10'b0111101001;
  /* fppowtf32.vhdl:1608:24  */
  assign n5835 = x == 10'b0111101010;
  /* fppowtf32.vhdl:1609:24  */
  assign n5838 = x == 10'b0111101011;
  /* fppowtf32.vhdl:1610:24  */
  assign n5841 = x == 10'b0111101100;
  /* fppowtf32.vhdl:1611:24  */
  assign n5844 = x == 10'b0111101101;
  /* fppowtf32.vhdl:1612:24  */
  assign n5847 = x == 10'b0111101110;
  /* fppowtf32.vhdl:1613:24  */
  assign n5850 = x == 10'b0111101111;
  /* fppowtf32.vhdl:1614:24  */
  assign n5853 = x == 10'b0111110000;
  /* fppowtf32.vhdl:1615:24  */
  assign n5856 = x == 10'b0111110001;
  /* fppowtf32.vhdl:1616:24  */
  assign n5859 = x == 10'b0111110010;
  /* fppowtf32.vhdl:1617:24  */
  assign n5862 = x == 10'b0111110011;
  /* fppowtf32.vhdl:1618:24  */
  assign n5865 = x == 10'b0111110100;
  /* fppowtf32.vhdl:1619:24  */
  assign n5868 = x == 10'b0111110101;
  /* fppowtf32.vhdl:1620:24  */
  assign n5871 = x == 10'b0111110110;
  /* fppowtf32.vhdl:1621:24  */
  assign n5874 = x == 10'b0111110111;
  /* fppowtf32.vhdl:1622:24  */
  assign n5877 = x == 10'b0111111000;
  /* fppowtf32.vhdl:1623:24  */
  assign n5880 = x == 10'b0111111001;
  /* fppowtf32.vhdl:1624:24  */
  assign n5883 = x == 10'b0111111010;
  /* fppowtf32.vhdl:1625:24  */
  assign n5886 = x == 10'b0111111011;
  /* fppowtf32.vhdl:1626:24  */
  assign n5889 = x == 10'b0111111100;
  /* fppowtf32.vhdl:1627:24  */
  assign n5892 = x == 10'b0111111101;
  /* fppowtf32.vhdl:1628:24  */
  assign n5895 = x == 10'b0111111110;
  /* fppowtf32.vhdl:1629:24  */
  assign n5898 = x == 10'b0111111111;
  /* fppowtf32.vhdl:1630:24  */
  assign n5901 = x == 10'b1000000000;
  /* fppowtf32.vhdl:1631:24  */
  assign n5904 = x == 10'b1000000001;
  /* fppowtf32.vhdl:1632:24  */
  assign n5907 = x == 10'b1000000010;
  /* fppowtf32.vhdl:1633:24  */
  assign n5910 = x == 10'b1000000011;
  /* fppowtf32.vhdl:1634:24  */
  assign n5913 = x == 10'b1000000100;
  /* fppowtf32.vhdl:1635:24  */
  assign n5916 = x == 10'b1000000101;
  /* fppowtf32.vhdl:1636:24  */
  assign n5919 = x == 10'b1000000110;
  /* fppowtf32.vhdl:1637:24  */
  assign n5922 = x == 10'b1000000111;
  /* fppowtf32.vhdl:1638:24  */
  assign n5925 = x == 10'b1000001000;
  /* fppowtf32.vhdl:1639:24  */
  assign n5928 = x == 10'b1000001001;
  /* fppowtf32.vhdl:1640:24  */
  assign n5931 = x == 10'b1000001010;
  /* fppowtf32.vhdl:1641:24  */
  assign n5934 = x == 10'b1000001011;
  /* fppowtf32.vhdl:1642:24  */
  assign n5937 = x == 10'b1000001100;
  /* fppowtf32.vhdl:1643:24  */
  assign n5940 = x == 10'b1000001101;
  /* fppowtf32.vhdl:1644:24  */
  assign n5943 = x == 10'b1000001110;
  /* fppowtf32.vhdl:1645:24  */
  assign n5946 = x == 10'b1000001111;
  /* fppowtf32.vhdl:1646:24  */
  assign n5949 = x == 10'b1000010000;
  /* fppowtf32.vhdl:1647:24  */
  assign n5952 = x == 10'b1000010001;
  /* fppowtf32.vhdl:1648:24  */
  assign n5955 = x == 10'b1000010010;
  /* fppowtf32.vhdl:1649:24  */
  assign n5958 = x == 10'b1000010011;
  /* fppowtf32.vhdl:1650:24  */
  assign n5961 = x == 10'b1000010100;
  /* fppowtf32.vhdl:1651:24  */
  assign n5964 = x == 10'b1000010101;
  /* fppowtf32.vhdl:1652:24  */
  assign n5967 = x == 10'b1000010110;
  /* fppowtf32.vhdl:1653:24  */
  assign n5970 = x == 10'b1000010111;
  /* fppowtf32.vhdl:1654:24  */
  assign n5973 = x == 10'b1000011000;
  /* fppowtf32.vhdl:1655:24  */
  assign n5976 = x == 10'b1000011001;
  /* fppowtf32.vhdl:1656:24  */
  assign n5979 = x == 10'b1000011010;
  /* fppowtf32.vhdl:1657:24  */
  assign n5982 = x == 10'b1000011011;
  /* fppowtf32.vhdl:1658:24  */
  assign n5985 = x == 10'b1000011100;
  /* fppowtf32.vhdl:1659:24  */
  assign n5988 = x == 10'b1000011101;
  /* fppowtf32.vhdl:1660:24  */
  assign n5991 = x == 10'b1000011110;
  /* fppowtf32.vhdl:1661:24  */
  assign n5994 = x == 10'b1000011111;
  /* fppowtf32.vhdl:1662:24  */
  assign n5997 = x == 10'b1000100000;
  /* fppowtf32.vhdl:1663:24  */
  assign n6000 = x == 10'b1000100001;
  /* fppowtf32.vhdl:1664:24  */
  assign n6003 = x == 10'b1000100010;
  /* fppowtf32.vhdl:1665:24  */
  assign n6006 = x == 10'b1000100011;
  /* fppowtf32.vhdl:1666:24  */
  assign n6009 = x == 10'b1000100100;
  /* fppowtf32.vhdl:1667:24  */
  assign n6012 = x == 10'b1000100101;
  /* fppowtf32.vhdl:1668:24  */
  assign n6015 = x == 10'b1000100110;
  /* fppowtf32.vhdl:1669:24  */
  assign n6018 = x == 10'b1000100111;
  /* fppowtf32.vhdl:1670:24  */
  assign n6021 = x == 10'b1000101000;
  /* fppowtf32.vhdl:1671:24  */
  assign n6024 = x == 10'b1000101001;
  /* fppowtf32.vhdl:1672:24  */
  assign n6027 = x == 10'b1000101010;
  /* fppowtf32.vhdl:1673:24  */
  assign n6030 = x == 10'b1000101011;
  /* fppowtf32.vhdl:1674:24  */
  assign n6033 = x == 10'b1000101100;
  /* fppowtf32.vhdl:1675:24  */
  assign n6036 = x == 10'b1000101101;
  /* fppowtf32.vhdl:1676:24  */
  assign n6039 = x == 10'b1000101110;
  /* fppowtf32.vhdl:1677:24  */
  assign n6042 = x == 10'b1000101111;
  /* fppowtf32.vhdl:1678:24  */
  assign n6045 = x == 10'b1000110000;
  /* fppowtf32.vhdl:1679:24  */
  assign n6048 = x == 10'b1000110001;
  /* fppowtf32.vhdl:1680:24  */
  assign n6051 = x == 10'b1000110010;
  /* fppowtf32.vhdl:1681:24  */
  assign n6054 = x == 10'b1000110011;
  /* fppowtf32.vhdl:1682:24  */
  assign n6057 = x == 10'b1000110100;
  /* fppowtf32.vhdl:1683:24  */
  assign n6060 = x == 10'b1000110101;
  /* fppowtf32.vhdl:1684:24  */
  assign n6063 = x == 10'b1000110110;
  /* fppowtf32.vhdl:1685:24  */
  assign n6066 = x == 10'b1000110111;
  /* fppowtf32.vhdl:1686:24  */
  assign n6069 = x == 10'b1000111000;
  /* fppowtf32.vhdl:1687:24  */
  assign n6072 = x == 10'b1000111001;
  /* fppowtf32.vhdl:1688:24  */
  assign n6075 = x == 10'b1000111010;
  /* fppowtf32.vhdl:1689:24  */
  assign n6078 = x == 10'b1000111011;
  /* fppowtf32.vhdl:1690:24  */
  assign n6081 = x == 10'b1000111100;
  /* fppowtf32.vhdl:1691:24  */
  assign n6084 = x == 10'b1000111101;
  /* fppowtf32.vhdl:1692:24  */
  assign n6087 = x == 10'b1000111110;
  /* fppowtf32.vhdl:1693:24  */
  assign n6090 = x == 10'b1000111111;
  /* fppowtf32.vhdl:1694:24  */
  assign n6093 = x == 10'b1001000000;
  /* fppowtf32.vhdl:1695:24  */
  assign n6096 = x == 10'b1001000001;
  /* fppowtf32.vhdl:1696:24  */
  assign n6099 = x == 10'b1001000010;
  /* fppowtf32.vhdl:1697:24  */
  assign n6102 = x == 10'b1001000011;
  /* fppowtf32.vhdl:1698:24  */
  assign n6105 = x == 10'b1001000100;
  /* fppowtf32.vhdl:1699:24  */
  assign n6108 = x == 10'b1001000101;
  /* fppowtf32.vhdl:1700:24  */
  assign n6111 = x == 10'b1001000110;
  /* fppowtf32.vhdl:1701:24  */
  assign n6114 = x == 10'b1001000111;
  /* fppowtf32.vhdl:1702:24  */
  assign n6117 = x == 10'b1001001000;
  /* fppowtf32.vhdl:1703:24  */
  assign n6120 = x == 10'b1001001001;
  /* fppowtf32.vhdl:1704:24  */
  assign n6123 = x == 10'b1001001010;
  /* fppowtf32.vhdl:1705:24  */
  assign n6126 = x == 10'b1001001011;
  /* fppowtf32.vhdl:1706:24  */
  assign n6129 = x == 10'b1001001100;
  /* fppowtf32.vhdl:1707:24  */
  assign n6132 = x == 10'b1001001101;
  /* fppowtf32.vhdl:1708:24  */
  assign n6135 = x == 10'b1001001110;
  /* fppowtf32.vhdl:1709:24  */
  assign n6138 = x == 10'b1001001111;
  /* fppowtf32.vhdl:1710:24  */
  assign n6141 = x == 10'b1001010000;
  /* fppowtf32.vhdl:1711:24  */
  assign n6144 = x == 10'b1001010001;
  /* fppowtf32.vhdl:1712:24  */
  assign n6147 = x == 10'b1001010010;
  /* fppowtf32.vhdl:1713:24  */
  assign n6150 = x == 10'b1001010011;
  /* fppowtf32.vhdl:1714:24  */
  assign n6153 = x == 10'b1001010100;
  /* fppowtf32.vhdl:1715:24  */
  assign n6156 = x == 10'b1001010101;
  /* fppowtf32.vhdl:1716:24  */
  assign n6159 = x == 10'b1001010110;
  /* fppowtf32.vhdl:1717:24  */
  assign n6162 = x == 10'b1001010111;
  /* fppowtf32.vhdl:1718:24  */
  assign n6165 = x == 10'b1001011000;
  /* fppowtf32.vhdl:1719:24  */
  assign n6168 = x == 10'b1001011001;
  /* fppowtf32.vhdl:1720:24  */
  assign n6171 = x == 10'b1001011010;
  /* fppowtf32.vhdl:1721:24  */
  assign n6174 = x == 10'b1001011011;
  /* fppowtf32.vhdl:1722:24  */
  assign n6177 = x == 10'b1001011100;
  /* fppowtf32.vhdl:1723:24  */
  assign n6180 = x == 10'b1001011101;
  /* fppowtf32.vhdl:1724:24  */
  assign n6183 = x == 10'b1001011110;
  /* fppowtf32.vhdl:1725:24  */
  assign n6186 = x == 10'b1001011111;
  /* fppowtf32.vhdl:1726:24  */
  assign n6189 = x == 10'b1001100000;
  /* fppowtf32.vhdl:1727:24  */
  assign n6192 = x == 10'b1001100001;
  /* fppowtf32.vhdl:1728:24  */
  assign n6195 = x == 10'b1001100010;
  /* fppowtf32.vhdl:1729:24  */
  assign n6198 = x == 10'b1001100011;
  /* fppowtf32.vhdl:1730:24  */
  assign n6201 = x == 10'b1001100100;
  /* fppowtf32.vhdl:1731:24  */
  assign n6204 = x == 10'b1001100101;
  /* fppowtf32.vhdl:1732:24  */
  assign n6207 = x == 10'b1001100110;
  /* fppowtf32.vhdl:1733:24  */
  assign n6210 = x == 10'b1001100111;
  /* fppowtf32.vhdl:1734:24  */
  assign n6213 = x == 10'b1001101000;
  /* fppowtf32.vhdl:1735:24  */
  assign n6216 = x == 10'b1001101001;
  /* fppowtf32.vhdl:1736:24  */
  assign n6219 = x == 10'b1001101010;
  /* fppowtf32.vhdl:1737:24  */
  assign n6222 = x == 10'b1001101011;
  /* fppowtf32.vhdl:1738:24  */
  assign n6225 = x == 10'b1001101100;
  /* fppowtf32.vhdl:1739:24  */
  assign n6228 = x == 10'b1001101101;
  /* fppowtf32.vhdl:1740:24  */
  assign n6231 = x == 10'b1001101110;
  /* fppowtf32.vhdl:1741:24  */
  assign n6234 = x == 10'b1001101111;
  /* fppowtf32.vhdl:1742:24  */
  assign n6237 = x == 10'b1001110000;
  /* fppowtf32.vhdl:1743:24  */
  assign n6240 = x == 10'b1001110001;
  /* fppowtf32.vhdl:1744:24  */
  assign n6243 = x == 10'b1001110010;
  /* fppowtf32.vhdl:1745:24  */
  assign n6246 = x == 10'b1001110011;
  /* fppowtf32.vhdl:1746:24  */
  assign n6249 = x == 10'b1001110100;
  /* fppowtf32.vhdl:1747:24  */
  assign n6252 = x == 10'b1001110101;
  /* fppowtf32.vhdl:1748:24  */
  assign n6255 = x == 10'b1001110110;
  /* fppowtf32.vhdl:1749:24  */
  assign n6258 = x == 10'b1001110111;
  /* fppowtf32.vhdl:1750:24  */
  assign n6261 = x == 10'b1001111000;
  /* fppowtf32.vhdl:1751:24  */
  assign n6264 = x == 10'b1001111001;
  /* fppowtf32.vhdl:1752:24  */
  assign n6267 = x == 10'b1001111010;
  /* fppowtf32.vhdl:1753:24  */
  assign n6270 = x == 10'b1001111011;
  /* fppowtf32.vhdl:1754:24  */
  assign n6273 = x == 10'b1001111100;
  /* fppowtf32.vhdl:1755:24  */
  assign n6276 = x == 10'b1001111101;
  /* fppowtf32.vhdl:1756:24  */
  assign n6279 = x == 10'b1001111110;
  /* fppowtf32.vhdl:1757:24  */
  assign n6282 = x == 10'b1001111111;
  /* fppowtf32.vhdl:1758:24  */
  assign n6285 = x == 10'b1010000000;
  /* fppowtf32.vhdl:1759:24  */
  assign n6288 = x == 10'b1010000001;
  /* fppowtf32.vhdl:1760:24  */
  assign n6291 = x == 10'b1010000010;
  /* fppowtf32.vhdl:1761:24  */
  assign n6294 = x == 10'b1010000011;
  /* fppowtf32.vhdl:1762:24  */
  assign n6297 = x == 10'b1010000100;
  /* fppowtf32.vhdl:1763:24  */
  assign n6300 = x == 10'b1010000101;
  /* fppowtf32.vhdl:1764:24  */
  assign n6303 = x == 10'b1010000110;
  /* fppowtf32.vhdl:1765:24  */
  assign n6306 = x == 10'b1010000111;
  /* fppowtf32.vhdl:1766:24  */
  assign n6309 = x == 10'b1010001000;
  /* fppowtf32.vhdl:1767:24  */
  assign n6312 = x == 10'b1010001001;
  /* fppowtf32.vhdl:1768:24  */
  assign n6315 = x == 10'b1010001010;
  /* fppowtf32.vhdl:1769:24  */
  assign n6318 = x == 10'b1010001011;
  /* fppowtf32.vhdl:1770:24  */
  assign n6321 = x == 10'b1010001100;
  /* fppowtf32.vhdl:1771:24  */
  assign n6324 = x == 10'b1010001101;
  /* fppowtf32.vhdl:1772:24  */
  assign n6327 = x == 10'b1010001110;
  /* fppowtf32.vhdl:1773:24  */
  assign n6330 = x == 10'b1010001111;
  /* fppowtf32.vhdl:1774:24  */
  assign n6333 = x == 10'b1010010000;
  /* fppowtf32.vhdl:1775:24  */
  assign n6336 = x == 10'b1010010001;
  /* fppowtf32.vhdl:1776:24  */
  assign n6339 = x == 10'b1010010010;
  /* fppowtf32.vhdl:1777:24  */
  assign n6342 = x == 10'b1010010011;
  /* fppowtf32.vhdl:1778:24  */
  assign n6345 = x == 10'b1010010100;
  /* fppowtf32.vhdl:1779:24  */
  assign n6348 = x == 10'b1010010101;
  /* fppowtf32.vhdl:1780:24  */
  assign n6351 = x == 10'b1010010110;
  /* fppowtf32.vhdl:1781:24  */
  assign n6354 = x == 10'b1010010111;
  /* fppowtf32.vhdl:1782:24  */
  assign n6357 = x == 10'b1010011000;
  /* fppowtf32.vhdl:1783:24  */
  assign n6360 = x == 10'b1010011001;
  /* fppowtf32.vhdl:1784:24  */
  assign n6363 = x == 10'b1010011010;
  /* fppowtf32.vhdl:1785:24  */
  assign n6366 = x == 10'b1010011011;
  /* fppowtf32.vhdl:1786:24  */
  assign n6369 = x == 10'b1010011100;
  /* fppowtf32.vhdl:1787:24  */
  assign n6372 = x == 10'b1010011101;
  /* fppowtf32.vhdl:1788:24  */
  assign n6375 = x == 10'b1010011110;
  /* fppowtf32.vhdl:1789:24  */
  assign n6378 = x == 10'b1010011111;
  /* fppowtf32.vhdl:1790:24  */
  assign n6381 = x == 10'b1010100000;
  /* fppowtf32.vhdl:1791:24  */
  assign n6384 = x == 10'b1010100001;
  /* fppowtf32.vhdl:1792:24  */
  assign n6387 = x == 10'b1010100010;
  /* fppowtf32.vhdl:1793:24  */
  assign n6390 = x == 10'b1010100011;
  /* fppowtf32.vhdl:1794:24  */
  assign n6393 = x == 10'b1010100100;
  /* fppowtf32.vhdl:1795:24  */
  assign n6396 = x == 10'b1010100101;
  /* fppowtf32.vhdl:1796:24  */
  assign n6399 = x == 10'b1010100110;
  /* fppowtf32.vhdl:1797:24  */
  assign n6402 = x == 10'b1010100111;
  /* fppowtf32.vhdl:1798:24  */
  assign n6405 = x == 10'b1010101000;
  /* fppowtf32.vhdl:1799:24  */
  assign n6408 = x == 10'b1010101001;
  /* fppowtf32.vhdl:1800:24  */
  assign n6411 = x == 10'b1010101010;
  /* fppowtf32.vhdl:1801:24  */
  assign n6414 = x == 10'b1010101011;
  /* fppowtf32.vhdl:1802:24  */
  assign n6417 = x == 10'b1010101100;
  /* fppowtf32.vhdl:1803:24  */
  assign n6420 = x == 10'b1010101101;
  /* fppowtf32.vhdl:1804:24  */
  assign n6423 = x == 10'b1010101110;
  /* fppowtf32.vhdl:1805:24  */
  assign n6426 = x == 10'b1010101111;
  /* fppowtf32.vhdl:1806:24  */
  assign n6429 = x == 10'b1010110000;
  /* fppowtf32.vhdl:1807:24  */
  assign n6432 = x == 10'b1010110001;
  /* fppowtf32.vhdl:1808:24  */
  assign n6435 = x == 10'b1010110010;
  /* fppowtf32.vhdl:1809:24  */
  assign n6438 = x == 10'b1010110011;
  /* fppowtf32.vhdl:1810:24  */
  assign n6441 = x == 10'b1010110100;
  /* fppowtf32.vhdl:1811:24  */
  assign n6444 = x == 10'b1010110101;
  /* fppowtf32.vhdl:1812:24  */
  assign n6447 = x == 10'b1010110110;
  /* fppowtf32.vhdl:1813:24  */
  assign n6450 = x == 10'b1010110111;
  /* fppowtf32.vhdl:1814:24  */
  assign n6453 = x == 10'b1010111000;
  /* fppowtf32.vhdl:1815:24  */
  assign n6456 = x == 10'b1010111001;
  /* fppowtf32.vhdl:1816:24  */
  assign n6459 = x == 10'b1010111010;
  /* fppowtf32.vhdl:1817:24  */
  assign n6462 = x == 10'b1010111011;
  /* fppowtf32.vhdl:1818:24  */
  assign n6465 = x == 10'b1010111100;
  /* fppowtf32.vhdl:1819:24  */
  assign n6468 = x == 10'b1010111101;
  /* fppowtf32.vhdl:1820:24  */
  assign n6471 = x == 10'b1010111110;
  /* fppowtf32.vhdl:1821:24  */
  assign n6474 = x == 10'b1010111111;
  /* fppowtf32.vhdl:1822:24  */
  assign n6477 = x == 10'b1011000000;
  /* fppowtf32.vhdl:1823:24  */
  assign n6480 = x == 10'b1011000001;
  /* fppowtf32.vhdl:1824:24  */
  assign n6483 = x == 10'b1011000010;
  /* fppowtf32.vhdl:1825:24  */
  assign n6486 = x == 10'b1011000011;
  /* fppowtf32.vhdl:1826:24  */
  assign n6489 = x == 10'b1011000100;
  /* fppowtf32.vhdl:1827:24  */
  assign n6492 = x == 10'b1011000101;
  /* fppowtf32.vhdl:1828:24  */
  assign n6495 = x == 10'b1011000110;
  /* fppowtf32.vhdl:1829:24  */
  assign n6498 = x == 10'b1011000111;
  /* fppowtf32.vhdl:1830:24  */
  assign n6501 = x == 10'b1011001000;
  /* fppowtf32.vhdl:1831:24  */
  assign n6504 = x == 10'b1011001001;
  /* fppowtf32.vhdl:1832:24  */
  assign n6507 = x == 10'b1011001010;
  /* fppowtf32.vhdl:1833:24  */
  assign n6510 = x == 10'b1011001011;
  /* fppowtf32.vhdl:1834:24  */
  assign n6513 = x == 10'b1011001100;
  /* fppowtf32.vhdl:1835:24  */
  assign n6516 = x == 10'b1011001101;
  /* fppowtf32.vhdl:1836:24  */
  assign n6519 = x == 10'b1011001110;
  /* fppowtf32.vhdl:1837:24  */
  assign n6522 = x == 10'b1011001111;
  /* fppowtf32.vhdl:1838:24  */
  assign n6525 = x == 10'b1011010000;
  /* fppowtf32.vhdl:1839:24  */
  assign n6528 = x == 10'b1011010001;
  /* fppowtf32.vhdl:1840:24  */
  assign n6531 = x == 10'b1011010010;
  /* fppowtf32.vhdl:1841:24  */
  assign n6534 = x == 10'b1011010011;
  /* fppowtf32.vhdl:1842:24  */
  assign n6537 = x == 10'b1011010100;
  /* fppowtf32.vhdl:1843:24  */
  assign n6540 = x == 10'b1011010101;
  /* fppowtf32.vhdl:1844:24  */
  assign n6543 = x == 10'b1011010110;
  /* fppowtf32.vhdl:1845:24  */
  assign n6546 = x == 10'b1011010111;
  /* fppowtf32.vhdl:1846:24  */
  assign n6549 = x == 10'b1011011000;
  /* fppowtf32.vhdl:1847:24  */
  assign n6552 = x == 10'b1011011001;
  /* fppowtf32.vhdl:1848:24  */
  assign n6555 = x == 10'b1011011010;
  /* fppowtf32.vhdl:1849:24  */
  assign n6558 = x == 10'b1011011011;
  /* fppowtf32.vhdl:1850:24  */
  assign n6561 = x == 10'b1011011100;
  /* fppowtf32.vhdl:1851:24  */
  assign n6564 = x == 10'b1011011101;
  /* fppowtf32.vhdl:1852:24  */
  assign n6567 = x == 10'b1011011110;
  /* fppowtf32.vhdl:1853:24  */
  assign n6570 = x == 10'b1011011111;
  /* fppowtf32.vhdl:1854:24  */
  assign n6573 = x == 10'b1011100000;
  /* fppowtf32.vhdl:1855:24  */
  assign n6576 = x == 10'b1011100001;
  /* fppowtf32.vhdl:1856:24  */
  assign n6579 = x == 10'b1011100010;
  /* fppowtf32.vhdl:1857:24  */
  assign n6582 = x == 10'b1011100011;
  /* fppowtf32.vhdl:1858:24  */
  assign n6585 = x == 10'b1011100100;
  /* fppowtf32.vhdl:1859:24  */
  assign n6588 = x == 10'b1011100101;
  /* fppowtf32.vhdl:1860:24  */
  assign n6591 = x == 10'b1011100110;
  /* fppowtf32.vhdl:1861:24  */
  assign n6594 = x == 10'b1011100111;
  /* fppowtf32.vhdl:1862:24  */
  assign n6597 = x == 10'b1011101000;
  /* fppowtf32.vhdl:1863:24  */
  assign n6600 = x == 10'b1011101001;
  /* fppowtf32.vhdl:1864:24  */
  assign n6603 = x == 10'b1011101010;
  /* fppowtf32.vhdl:1865:24  */
  assign n6606 = x == 10'b1011101011;
  /* fppowtf32.vhdl:1866:24  */
  assign n6609 = x == 10'b1011101100;
  /* fppowtf32.vhdl:1867:24  */
  assign n6612 = x == 10'b1011101101;
  /* fppowtf32.vhdl:1868:24  */
  assign n6615 = x == 10'b1011101110;
  /* fppowtf32.vhdl:1869:24  */
  assign n6618 = x == 10'b1011101111;
  /* fppowtf32.vhdl:1870:24  */
  assign n6621 = x == 10'b1011110000;
  /* fppowtf32.vhdl:1871:24  */
  assign n6624 = x == 10'b1011110001;
  /* fppowtf32.vhdl:1872:24  */
  assign n6627 = x == 10'b1011110010;
  /* fppowtf32.vhdl:1873:24  */
  assign n6630 = x == 10'b1011110011;
  /* fppowtf32.vhdl:1874:24  */
  assign n6633 = x == 10'b1011110100;
  /* fppowtf32.vhdl:1875:24  */
  assign n6636 = x == 10'b1011110101;
  /* fppowtf32.vhdl:1876:24  */
  assign n6639 = x == 10'b1011110110;
  /* fppowtf32.vhdl:1877:24  */
  assign n6642 = x == 10'b1011110111;
  /* fppowtf32.vhdl:1878:24  */
  assign n6645 = x == 10'b1011111000;
  /* fppowtf32.vhdl:1879:24  */
  assign n6648 = x == 10'b1011111001;
  /* fppowtf32.vhdl:1880:24  */
  assign n6651 = x == 10'b1011111010;
  /* fppowtf32.vhdl:1881:24  */
  assign n6654 = x == 10'b1011111011;
  /* fppowtf32.vhdl:1882:24  */
  assign n6657 = x == 10'b1011111100;
  /* fppowtf32.vhdl:1883:24  */
  assign n6660 = x == 10'b1011111101;
  /* fppowtf32.vhdl:1884:24  */
  assign n6663 = x == 10'b1011111110;
  /* fppowtf32.vhdl:1885:24  */
  assign n6666 = x == 10'b1011111111;
  /* fppowtf32.vhdl:1886:24  */
  assign n6669 = x == 10'b1100000000;
  /* fppowtf32.vhdl:1887:24  */
  assign n6672 = x == 10'b1100000001;
  /* fppowtf32.vhdl:1888:24  */
  assign n6675 = x == 10'b1100000010;
  /* fppowtf32.vhdl:1889:24  */
  assign n6678 = x == 10'b1100000011;
  /* fppowtf32.vhdl:1890:24  */
  assign n6681 = x == 10'b1100000100;
  /* fppowtf32.vhdl:1891:24  */
  assign n6684 = x == 10'b1100000101;
  /* fppowtf32.vhdl:1892:24  */
  assign n6687 = x == 10'b1100000110;
  /* fppowtf32.vhdl:1893:24  */
  assign n6690 = x == 10'b1100000111;
  /* fppowtf32.vhdl:1894:24  */
  assign n6693 = x == 10'b1100001000;
  /* fppowtf32.vhdl:1895:24  */
  assign n6696 = x == 10'b1100001001;
  /* fppowtf32.vhdl:1896:24  */
  assign n6699 = x == 10'b1100001010;
  /* fppowtf32.vhdl:1897:24  */
  assign n6702 = x == 10'b1100001011;
  /* fppowtf32.vhdl:1898:24  */
  assign n6705 = x == 10'b1100001100;
  /* fppowtf32.vhdl:1899:24  */
  assign n6708 = x == 10'b1100001101;
  /* fppowtf32.vhdl:1900:24  */
  assign n6711 = x == 10'b1100001110;
  /* fppowtf32.vhdl:1901:24  */
  assign n6714 = x == 10'b1100001111;
  /* fppowtf32.vhdl:1902:24  */
  assign n6717 = x == 10'b1100010000;
  /* fppowtf32.vhdl:1903:24  */
  assign n6720 = x == 10'b1100010001;
  /* fppowtf32.vhdl:1904:24  */
  assign n6723 = x == 10'b1100010010;
  /* fppowtf32.vhdl:1905:24  */
  assign n6726 = x == 10'b1100010011;
  /* fppowtf32.vhdl:1906:24  */
  assign n6729 = x == 10'b1100010100;
  /* fppowtf32.vhdl:1907:24  */
  assign n6732 = x == 10'b1100010101;
  /* fppowtf32.vhdl:1908:24  */
  assign n6735 = x == 10'b1100010110;
  /* fppowtf32.vhdl:1909:24  */
  assign n6738 = x == 10'b1100010111;
  /* fppowtf32.vhdl:1910:24  */
  assign n6741 = x == 10'b1100011000;
  /* fppowtf32.vhdl:1911:24  */
  assign n6744 = x == 10'b1100011001;
  /* fppowtf32.vhdl:1912:24  */
  assign n6747 = x == 10'b1100011010;
  /* fppowtf32.vhdl:1913:24  */
  assign n6750 = x == 10'b1100011011;
  /* fppowtf32.vhdl:1914:24  */
  assign n6753 = x == 10'b1100011100;
  /* fppowtf32.vhdl:1915:24  */
  assign n6756 = x == 10'b1100011101;
  /* fppowtf32.vhdl:1916:24  */
  assign n6759 = x == 10'b1100011110;
  /* fppowtf32.vhdl:1917:24  */
  assign n6762 = x == 10'b1100011111;
  /* fppowtf32.vhdl:1918:24  */
  assign n6765 = x == 10'b1100100000;
  /* fppowtf32.vhdl:1919:24  */
  assign n6768 = x == 10'b1100100001;
  /* fppowtf32.vhdl:1920:24  */
  assign n6771 = x == 10'b1100100010;
  /* fppowtf32.vhdl:1921:24  */
  assign n6774 = x == 10'b1100100011;
  /* fppowtf32.vhdl:1922:24  */
  assign n6777 = x == 10'b1100100100;
  /* fppowtf32.vhdl:1923:24  */
  assign n6780 = x == 10'b1100100101;
  /* fppowtf32.vhdl:1924:24  */
  assign n6783 = x == 10'b1100100110;
  /* fppowtf32.vhdl:1925:24  */
  assign n6786 = x == 10'b1100100111;
  /* fppowtf32.vhdl:1926:24  */
  assign n6789 = x == 10'b1100101000;
  /* fppowtf32.vhdl:1927:24  */
  assign n6792 = x == 10'b1100101001;
  /* fppowtf32.vhdl:1928:24  */
  assign n6795 = x == 10'b1100101010;
  /* fppowtf32.vhdl:1929:24  */
  assign n6798 = x == 10'b1100101011;
  /* fppowtf32.vhdl:1930:24  */
  assign n6801 = x == 10'b1100101100;
  /* fppowtf32.vhdl:1931:24  */
  assign n6804 = x == 10'b1100101101;
  /* fppowtf32.vhdl:1932:24  */
  assign n6807 = x == 10'b1100101110;
  /* fppowtf32.vhdl:1933:24  */
  assign n6810 = x == 10'b1100101111;
  /* fppowtf32.vhdl:1934:24  */
  assign n6813 = x == 10'b1100110000;
  /* fppowtf32.vhdl:1935:24  */
  assign n6816 = x == 10'b1100110001;
  /* fppowtf32.vhdl:1936:24  */
  assign n6819 = x == 10'b1100110010;
  /* fppowtf32.vhdl:1937:24  */
  assign n6822 = x == 10'b1100110011;
  /* fppowtf32.vhdl:1938:24  */
  assign n6825 = x == 10'b1100110100;
  /* fppowtf32.vhdl:1939:24  */
  assign n6828 = x == 10'b1100110101;
  /* fppowtf32.vhdl:1940:24  */
  assign n6831 = x == 10'b1100110110;
  /* fppowtf32.vhdl:1941:24  */
  assign n6834 = x == 10'b1100110111;
  /* fppowtf32.vhdl:1942:24  */
  assign n6837 = x == 10'b1100111000;
  /* fppowtf32.vhdl:1943:24  */
  assign n6840 = x == 10'b1100111001;
  /* fppowtf32.vhdl:1944:24  */
  assign n6843 = x == 10'b1100111010;
  /* fppowtf32.vhdl:1945:24  */
  assign n6846 = x == 10'b1100111011;
  /* fppowtf32.vhdl:1946:24  */
  assign n6849 = x == 10'b1100111100;
  /* fppowtf32.vhdl:1947:24  */
  assign n6852 = x == 10'b1100111101;
  /* fppowtf32.vhdl:1948:24  */
  assign n6855 = x == 10'b1100111110;
  /* fppowtf32.vhdl:1949:24  */
  assign n6858 = x == 10'b1100111111;
  /* fppowtf32.vhdl:1950:24  */
  assign n6861 = x == 10'b1101000000;
  /* fppowtf32.vhdl:1951:24  */
  assign n6864 = x == 10'b1101000001;
  /* fppowtf32.vhdl:1952:24  */
  assign n6867 = x == 10'b1101000010;
  /* fppowtf32.vhdl:1953:24  */
  assign n6870 = x == 10'b1101000011;
  /* fppowtf32.vhdl:1954:24  */
  assign n6873 = x == 10'b1101000100;
  /* fppowtf32.vhdl:1955:24  */
  assign n6876 = x == 10'b1101000101;
  /* fppowtf32.vhdl:1956:24  */
  assign n6879 = x == 10'b1101000110;
  /* fppowtf32.vhdl:1957:24  */
  assign n6882 = x == 10'b1101000111;
  /* fppowtf32.vhdl:1958:24  */
  assign n6885 = x == 10'b1101001000;
  /* fppowtf32.vhdl:1959:24  */
  assign n6888 = x == 10'b1101001001;
  /* fppowtf32.vhdl:1960:24  */
  assign n6891 = x == 10'b1101001010;
  /* fppowtf32.vhdl:1961:24  */
  assign n6894 = x == 10'b1101001011;
  /* fppowtf32.vhdl:1962:24  */
  assign n6897 = x == 10'b1101001100;
  /* fppowtf32.vhdl:1963:24  */
  assign n6900 = x == 10'b1101001101;
  /* fppowtf32.vhdl:1964:24  */
  assign n6903 = x == 10'b1101001110;
  /* fppowtf32.vhdl:1965:24  */
  assign n6906 = x == 10'b1101001111;
  /* fppowtf32.vhdl:1966:24  */
  assign n6909 = x == 10'b1101010000;
  /* fppowtf32.vhdl:1967:24  */
  assign n6912 = x == 10'b1101010001;
  /* fppowtf32.vhdl:1968:24  */
  assign n6915 = x == 10'b1101010010;
  /* fppowtf32.vhdl:1969:24  */
  assign n6918 = x == 10'b1101010011;
  /* fppowtf32.vhdl:1970:24  */
  assign n6921 = x == 10'b1101010100;
  /* fppowtf32.vhdl:1971:24  */
  assign n6924 = x == 10'b1101010101;
  /* fppowtf32.vhdl:1972:24  */
  assign n6927 = x == 10'b1101010110;
  /* fppowtf32.vhdl:1973:24  */
  assign n6930 = x == 10'b1101010111;
  /* fppowtf32.vhdl:1974:24  */
  assign n6933 = x == 10'b1101011000;
  /* fppowtf32.vhdl:1975:24  */
  assign n6936 = x == 10'b1101011001;
  /* fppowtf32.vhdl:1976:24  */
  assign n6939 = x == 10'b1101011010;
  /* fppowtf32.vhdl:1977:24  */
  assign n6942 = x == 10'b1101011011;
  /* fppowtf32.vhdl:1978:24  */
  assign n6945 = x == 10'b1101011100;
  /* fppowtf32.vhdl:1979:24  */
  assign n6948 = x == 10'b1101011101;
  /* fppowtf32.vhdl:1980:24  */
  assign n6951 = x == 10'b1101011110;
  /* fppowtf32.vhdl:1981:24  */
  assign n6954 = x == 10'b1101011111;
  /* fppowtf32.vhdl:1982:24  */
  assign n6957 = x == 10'b1101100000;
  /* fppowtf32.vhdl:1983:24  */
  assign n6960 = x == 10'b1101100001;
  /* fppowtf32.vhdl:1984:24  */
  assign n6963 = x == 10'b1101100010;
  /* fppowtf32.vhdl:1985:24  */
  assign n6966 = x == 10'b1101100011;
  /* fppowtf32.vhdl:1986:24  */
  assign n6969 = x == 10'b1101100100;
  /* fppowtf32.vhdl:1987:24  */
  assign n6972 = x == 10'b1101100101;
  /* fppowtf32.vhdl:1988:24  */
  assign n6975 = x == 10'b1101100110;
  /* fppowtf32.vhdl:1989:24  */
  assign n6978 = x == 10'b1101100111;
  /* fppowtf32.vhdl:1990:24  */
  assign n6981 = x == 10'b1101101000;
  /* fppowtf32.vhdl:1991:24  */
  assign n6984 = x == 10'b1101101001;
  /* fppowtf32.vhdl:1992:24  */
  assign n6987 = x == 10'b1101101010;
  /* fppowtf32.vhdl:1993:24  */
  assign n6990 = x == 10'b1101101011;
  /* fppowtf32.vhdl:1994:24  */
  assign n6993 = x == 10'b1101101100;
  /* fppowtf32.vhdl:1995:24  */
  assign n6996 = x == 10'b1101101101;
  /* fppowtf32.vhdl:1996:24  */
  assign n6999 = x == 10'b1101101110;
  /* fppowtf32.vhdl:1997:24  */
  assign n7002 = x == 10'b1101101111;
  /* fppowtf32.vhdl:1998:24  */
  assign n7005 = x == 10'b1101110000;
  /* fppowtf32.vhdl:1999:24  */
  assign n7008 = x == 10'b1101110001;
  /* fppowtf32.vhdl:2000:24  */
  assign n7011 = x == 10'b1101110010;
  /* fppowtf32.vhdl:2001:24  */
  assign n7014 = x == 10'b1101110011;
  /* fppowtf32.vhdl:2002:24  */
  assign n7017 = x == 10'b1101110100;
  /* fppowtf32.vhdl:2003:24  */
  assign n7020 = x == 10'b1101110101;
  /* fppowtf32.vhdl:2004:24  */
  assign n7023 = x == 10'b1101110110;
  /* fppowtf32.vhdl:2005:24  */
  assign n7026 = x == 10'b1101110111;
  /* fppowtf32.vhdl:2006:24  */
  assign n7029 = x == 10'b1101111000;
  /* fppowtf32.vhdl:2007:24  */
  assign n7032 = x == 10'b1101111001;
  /* fppowtf32.vhdl:2008:24  */
  assign n7035 = x == 10'b1101111010;
  /* fppowtf32.vhdl:2009:24  */
  assign n7038 = x == 10'b1101111011;
  /* fppowtf32.vhdl:2010:24  */
  assign n7041 = x == 10'b1101111100;
  /* fppowtf32.vhdl:2011:24  */
  assign n7044 = x == 10'b1101111101;
  /* fppowtf32.vhdl:2012:24  */
  assign n7047 = x == 10'b1101111110;
  /* fppowtf32.vhdl:2013:24  */
  assign n7050 = x == 10'b1101111111;
  /* fppowtf32.vhdl:2014:24  */
  assign n7053 = x == 10'b1110000000;
  /* fppowtf32.vhdl:2015:24  */
  assign n7056 = x == 10'b1110000001;
  /* fppowtf32.vhdl:2016:24  */
  assign n7059 = x == 10'b1110000010;
  /* fppowtf32.vhdl:2017:24  */
  assign n7062 = x == 10'b1110000011;
  /* fppowtf32.vhdl:2018:24  */
  assign n7065 = x == 10'b1110000100;
  /* fppowtf32.vhdl:2019:24  */
  assign n7068 = x == 10'b1110000101;
  /* fppowtf32.vhdl:2020:24  */
  assign n7071 = x == 10'b1110000110;
  /* fppowtf32.vhdl:2021:24  */
  assign n7074 = x == 10'b1110000111;
  /* fppowtf32.vhdl:2022:24  */
  assign n7077 = x == 10'b1110001000;
  /* fppowtf32.vhdl:2023:24  */
  assign n7080 = x == 10'b1110001001;
  /* fppowtf32.vhdl:2024:24  */
  assign n7083 = x == 10'b1110001010;
  /* fppowtf32.vhdl:2025:24  */
  assign n7086 = x == 10'b1110001011;
  /* fppowtf32.vhdl:2026:24  */
  assign n7089 = x == 10'b1110001100;
  /* fppowtf32.vhdl:2027:24  */
  assign n7092 = x == 10'b1110001101;
  /* fppowtf32.vhdl:2028:24  */
  assign n7095 = x == 10'b1110001110;
  /* fppowtf32.vhdl:2029:24  */
  assign n7098 = x == 10'b1110001111;
  /* fppowtf32.vhdl:2030:24  */
  assign n7101 = x == 10'b1110010000;
  /* fppowtf32.vhdl:2031:24  */
  assign n7104 = x == 10'b1110010001;
  /* fppowtf32.vhdl:2032:24  */
  assign n7107 = x == 10'b1110010010;
  /* fppowtf32.vhdl:2033:24  */
  assign n7110 = x == 10'b1110010011;
  /* fppowtf32.vhdl:2034:24  */
  assign n7113 = x == 10'b1110010100;
  /* fppowtf32.vhdl:2035:24  */
  assign n7116 = x == 10'b1110010101;
  /* fppowtf32.vhdl:2036:24  */
  assign n7119 = x == 10'b1110010110;
  /* fppowtf32.vhdl:2037:24  */
  assign n7122 = x == 10'b1110010111;
  /* fppowtf32.vhdl:2038:24  */
  assign n7125 = x == 10'b1110011000;
  /* fppowtf32.vhdl:2039:24  */
  assign n7128 = x == 10'b1110011001;
  /* fppowtf32.vhdl:2040:24  */
  assign n7131 = x == 10'b1110011010;
  /* fppowtf32.vhdl:2041:24  */
  assign n7134 = x == 10'b1110011011;
  /* fppowtf32.vhdl:2042:24  */
  assign n7137 = x == 10'b1110011100;
  /* fppowtf32.vhdl:2043:24  */
  assign n7140 = x == 10'b1110011101;
  /* fppowtf32.vhdl:2044:24  */
  assign n7143 = x == 10'b1110011110;
  /* fppowtf32.vhdl:2045:24  */
  assign n7146 = x == 10'b1110011111;
  /* fppowtf32.vhdl:2046:24  */
  assign n7149 = x == 10'b1110100000;
  /* fppowtf32.vhdl:2047:24  */
  assign n7152 = x == 10'b1110100001;
  /* fppowtf32.vhdl:2048:24  */
  assign n7155 = x == 10'b1110100010;
  /* fppowtf32.vhdl:2049:24  */
  assign n7158 = x == 10'b1110100011;
  /* fppowtf32.vhdl:2050:24  */
  assign n7161 = x == 10'b1110100100;
  /* fppowtf32.vhdl:2051:24  */
  assign n7164 = x == 10'b1110100101;
  /* fppowtf32.vhdl:2052:24  */
  assign n7167 = x == 10'b1110100110;
  /* fppowtf32.vhdl:2053:24  */
  assign n7170 = x == 10'b1110100111;
  /* fppowtf32.vhdl:2054:24  */
  assign n7173 = x == 10'b1110101000;
  /* fppowtf32.vhdl:2055:24  */
  assign n7176 = x == 10'b1110101001;
  /* fppowtf32.vhdl:2056:24  */
  assign n7179 = x == 10'b1110101010;
  /* fppowtf32.vhdl:2057:24  */
  assign n7182 = x == 10'b1110101011;
  /* fppowtf32.vhdl:2058:24  */
  assign n7185 = x == 10'b1110101100;
  /* fppowtf32.vhdl:2059:24  */
  assign n7188 = x == 10'b1110101101;
  /* fppowtf32.vhdl:2060:24  */
  assign n7191 = x == 10'b1110101110;
  /* fppowtf32.vhdl:2061:24  */
  assign n7194 = x == 10'b1110101111;
  /* fppowtf32.vhdl:2062:24  */
  assign n7197 = x == 10'b1110110000;
  /* fppowtf32.vhdl:2063:24  */
  assign n7200 = x == 10'b1110110001;
  /* fppowtf32.vhdl:2064:24  */
  assign n7203 = x == 10'b1110110010;
  /* fppowtf32.vhdl:2065:24  */
  assign n7206 = x == 10'b1110110011;
  /* fppowtf32.vhdl:2066:24  */
  assign n7209 = x == 10'b1110110100;
  /* fppowtf32.vhdl:2067:24  */
  assign n7212 = x == 10'b1110110101;
  /* fppowtf32.vhdl:2068:24  */
  assign n7215 = x == 10'b1110110110;
  /* fppowtf32.vhdl:2069:24  */
  assign n7218 = x == 10'b1110110111;
  /* fppowtf32.vhdl:2070:24  */
  assign n7221 = x == 10'b1110111000;
  /* fppowtf32.vhdl:2071:24  */
  assign n7224 = x == 10'b1110111001;
  /* fppowtf32.vhdl:2072:24  */
  assign n7227 = x == 10'b1110111010;
  /* fppowtf32.vhdl:2073:24  */
  assign n7230 = x == 10'b1110111011;
  /* fppowtf32.vhdl:2074:24  */
  assign n7233 = x == 10'b1110111100;
  /* fppowtf32.vhdl:2075:24  */
  assign n7236 = x == 10'b1110111101;
  /* fppowtf32.vhdl:2076:24  */
  assign n7239 = x == 10'b1110111110;
  /* fppowtf32.vhdl:2077:24  */
  assign n7242 = x == 10'b1110111111;
  /* fppowtf32.vhdl:2078:24  */
  assign n7245 = x == 10'b1111000000;
  /* fppowtf32.vhdl:2079:24  */
  assign n7248 = x == 10'b1111000001;
  /* fppowtf32.vhdl:2080:24  */
  assign n7251 = x == 10'b1111000010;
  /* fppowtf32.vhdl:2081:24  */
  assign n7254 = x == 10'b1111000011;
  /* fppowtf32.vhdl:2082:24  */
  assign n7257 = x == 10'b1111000100;
  /* fppowtf32.vhdl:2083:24  */
  assign n7260 = x == 10'b1111000101;
  /* fppowtf32.vhdl:2084:24  */
  assign n7263 = x == 10'b1111000110;
  /* fppowtf32.vhdl:2085:24  */
  assign n7266 = x == 10'b1111000111;
  /* fppowtf32.vhdl:2086:24  */
  assign n7269 = x == 10'b1111001000;
  /* fppowtf32.vhdl:2087:24  */
  assign n7272 = x == 10'b1111001001;
  /* fppowtf32.vhdl:2088:24  */
  assign n7275 = x == 10'b1111001010;
  /* fppowtf32.vhdl:2089:24  */
  assign n7278 = x == 10'b1111001011;
  /* fppowtf32.vhdl:2090:24  */
  assign n7281 = x == 10'b1111001100;
  /* fppowtf32.vhdl:2091:24  */
  assign n7284 = x == 10'b1111001101;
  /* fppowtf32.vhdl:2092:24  */
  assign n7287 = x == 10'b1111001110;
  /* fppowtf32.vhdl:2093:24  */
  assign n7290 = x == 10'b1111001111;
  /* fppowtf32.vhdl:2094:24  */
  assign n7293 = x == 10'b1111010000;
  /* fppowtf32.vhdl:2095:24  */
  assign n7296 = x == 10'b1111010001;
  /* fppowtf32.vhdl:2096:24  */
  assign n7299 = x == 10'b1111010010;
  /* fppowtf32.vhdl:2097:24  */
  assign n7302 = x == 10'b1111010011;
  /* fppowtf32.vhdl:2098:24  */
  assign n7305 = x == 10'b1111010100;
  /* fppowtf32.vhdl:2099:24  */
  assign n7308 = x == 10'b1111010101;
  /* fppowtf32.vhdl:2100:24  */
  assign n7311 = x == 10'b1111010110;
  /* fppowtf32.vhdl:2101:24  */
  assign n7314 = x == 10'b1111010111;
  /* fppowtf32.vhdl:2102:24  */
  assign n7317 = x == 10'b1111011000;
  /* fppowtf32.vhdl:2103:24  */
  assign n7320 = x == 10'b1111011001;
  /* fppowtf32.vhdl:2104:24  */
  assign n7323 = x == 10'b1111011010;
  /* fppowtf32.vhdl:2105:24  */
  assign n7326 = x == 10'b1111011011;
  /* fppowtf32.vhdl:2106:24  */
  assign n7329 = x == 10'b1111011100;
  /* fppowtf32.vhdl:2107:24  */
  assign n7332 = x == 10'b1111011101;
  /* fppowtf32.vhdl:2108:24  */
  assign n7335 = x == 10'b1111011110;
  /* fppowtf32.vhdl:2109:24  */
  assign n7338 = x == 10'b1111011111;
  /* fppowtf32.vhdl:2110:24  */
  assign n7341 = x == 10'b1111100000;
  /* fppowtf32.vhdl:2111:24  */
  assign n7344 = x == 10'b1111100001;
  /* fppowtf32.vhdl:2112:24  */
  assign n7347 = x == 10'b1111100010;
  /* fppowtf32.vhdl:2113:24  */
  assign n7350 = x == 10'b1111100011;
  /* fppowtf32.vhdl:2114:24  */
  assign n7353 = x == 10'b1111100100;
  /* fppowtf32.vhdl:2115:24  */
  assign n7356 = x == 10'b1111100101;
  /* fppowtf32.vhdl:2116:24  */
  assign n7359 = x == 10'b1111100110;
  /* fppowtf32.vhdl:2117:24  */
  assign n7362 = x == 10'b1111100111;
  /* fppowtf32.vhdl:2118:24  */
  assign n7365 = x == 10'b1111101000;
  /* fppowtf32.vhdl:2119:24  */
  assign n7368 = x == 10'b1111101001;
  /* fppowtf32.vhdl:2120:24  */
  assign n7371 = x == 10'b1111101010;
  /* fppowtf32.vhdl:2121:24  */
  assign n7374 = x == 10'b1111101011;
  /* fppowtf32.vhdl:2122:24  */
  assign n7377 = x == 10'b1111101100;
  /* fppowtf32.vhdl:2123:24  */
  assign n7380 = x == 10'b1111101101;
  /* fppowtf32.vhdl:2124:24  */
  assign n7383 = x == 10'b1111101110;
  /* fppowtf32.vhdl:2125:24  */
  assign n7386 = x == 10'b1111101111;
  /* fppowtf32.vhdl:2126:24  */
  assign n7389 = x == 10'b1111110000;
  /* fppowtf32.vhdl:2127:24  */
  assign n7392 = x == 10'b1111110001;
  /* fppowtf32.vhdl:2128:24  */
  assign n7395 = x == 10'b1111110010;
  /* fppowtf32.vhdl:2129:24  */
  assign n7398 = x == 10'b1111110011;
  /* fppowtf32.vhdl:2130:24  */
  assign n7401 = x == 10'b1111110100;
  /* fppowtf32.vhdl:2131:24  */
  assign n7404 = x == 10'b1111110101;
  /* fppowtf32.vhdl:2132:24  */
  assign n7407 = x == 10'b1111110110;
  /* fppowtf32.vhdl:2133:24  */
  assign n7410 = x == 10'b1111110111;
  /* fppowtf32.vhdl:2134:24  */
  assign n7413 = x == 10'b1111111000;
  /* fppowtf32.vhdl:2135:24  */
  assign n7416 = x == 10'b1111111001;
  /* fppowtf32.vhdl:2136:24  */
  assign n7419 = x == 10'b1111111010;
  /* fppowtf32.vhdl:2137:24  */
  assign n7422 = x == 10'b1111111011;
  /* fppowtf32.vhdl:2138:24  */
  assign n7425 = x == 10'b1111111100;
  /* fppowtf32.vhdl:2139:24  */
  assign n7428 = x == 10'b1111111101;
  /* fppowtf32.vhdl:2140:24  */
  assign n7431 = x == 10'b1111111110;
  /* fppowtf32.vhdl:2141:24  */
  assign n7434 = x == 10'b1111111111;
  assign n7436 = {n7434, n7431, n7428, n7425, n7422, n7419, n7416, n7413, n7410, n7407, n7404, n7401, n7398, n7395, n7392, n7389, n7386, n7383, n7380, n7377, n7374, n7371, n7368, n7365, n7362, n7359, n7356, n7353, n7350, n7347, n7344, n7341, n7338, n7335, n7332, n7329, n7326, n7323, n7320, n7317, n7314, n7311, n7308, n7305, n7302, n7299, n7296, n7293, n7290, n7287, n7284, n7281, n7278, n7275, n7272, n7269, n7266, n7263, n7260, n7257, n7254, n7251, n7248, n7245, n7242, n7239, n7236, n7233, n7230, n7227, n7224, n7221, n7218, n7215, n7212, n7209, n7206, n7203, n7200, n7197, n7194, n7191, n7188, n7185, n7182, n7179, n7176, n7173, n7170, n7167, n7164, n7161, n7158, n7155, n7152, n7149, n7146, n7143, n7140, n7137, n7134, n7131, n7128, n7125, n7122, n7119, n7116, n7113, n7110, n7107, n7104, n7101, n7098, n7095, n7092, n7089, n7086, n7083, n7080, n7077, n7074, n7071, n7068, n7065, n7062, n7059, n7056, n7053, n7050, n7047, n7044, n7041, n7038, n7035, n7032, n7029, n7026, n7023, n7020, n7017, n7014, n7011, n7008, n7005, n7002, n6999, n6996, n6993, n6990, n6987, n6984, n6981, n6978, n6975, n6972, n6969, n6966, n6963, n6960, n6957, n6954, n6951, n6948, n6945, n6942, n6939, n6936, n6933, n6930, n6927, n6924, n6921, n6918, n6915, n6912, n6909, n6906, n6903, n6900, n6897, n6894, n6891, n6888, n6885, n6882, n6879, n6876, n6873, n6870, n6867, n6864, n6861, n6858, n6855, n6852, n6849, n6846, n6843, n6840, n6837, n6834, n6831, n6828, n6825, n6822, n6819, n6816, n6813, n6810, n6807, n6804, n6801, n6798, n6795, n6792, n6789, n6786, n6783, n6780, n6777, n6774, n6771, n6768, n6765, n6762, n6759, n6756, n6753, n6750, n6747, n6744, n6741, n6738, n6735, n6732, n6729, n6726, n6723, n6720, n6717, n6714, n6711, n6708, n6705, n6702, n6699, n6696, n6693, n6690, n6687, n6684, n6681, n6678, n6675, n6672, n6669, n6666, n6663, n6660, n6657, n6654, n6651, n6648, n6645, n6642, n6639, n6636, n6633, n6630, n6627, n6624, n6621, n6618, n6615, n6612, n6609, n6606, n6603, n6600, n6597, n6594, n6591, n6588, n6585, n6582, n6579, n6576, n6573, n6570, n6567, n6564, n6561, n6558, n6555, n6552, n6549, n6546, n6543, n6540, n6537, n6534, n6531, n6528, n6525, n6522, n6519, n6516, n6513, n6510, n6507, n6504, n6501, n6498, n6495, n6492, n6489, n6486, n6483, n6480, n6477, n6474, n6471, n6468, n6465, n6462, n6459, n6456, n6453, n6450, n6447, n6444, n6441, n6438, n6435, n6432, n6429, n6426, n6423, n6420, n6417, n6414, n6411, n6408, n6405, n6402, n6399, n6396, n6393, n6390, n6387, n6384, n6381, n6378, n6375, n6372, n6369, n6366, n6363, n6360, n6357, n6354, n6351, n6348, n6345, n6342, n6339, n6336, n6333, n6330, n6327, n6324, n6321, n6318, n6315, n6312, n6309, n6306, n6303, n6300, n6297, n6294, n6291, n6288, n6285, n6282, n6279, n6276, n6273, n6270, n6267, n6264, n6261, n6258, n6255, n6252, n6249, n6246, n6243, n6240, n6237, n6234, n6231, n6228, n6225, n6222, n6219, n6216, n6213, n6210, n6207, n6204, n6201, n6198, n6195, n6192, n6189, n6186, n6183, n6180, n6177, n6174, n6171, n6168, n6165, n6162, n6159, n6156, n6153, n6150, n6147, n6144, n6141, n6138, n6135, n6132, n6129, n6126, n6123, n6120, n6117, n6114, n6111, n6108, n6105, n6102, n6099, n6096, n6093, n6090, n6087, n6084, n6081, n6078, n6075, n6072, n6069, n6066, n6063, n6060, n6057, n6054, n6051, n6048, n6045, n6042, n6039, n6036, n6033, n6030, n6027, n6024, n6021, n6018, n6015, n6012, n6009, n6006, n6003, n6000, n5997, n5994, n5991, n5988, n5985, n5982, n5979, n5976, n5973, n5970, n5967, n5964, n5961, n5958, n5955, n5952, n5949, n5946, n5943, n5940, n5937, n5934, n5931, n5928, n5925, n5922, n5919, n5916, n5913, n5910, n5907, n5904, n5901, n5898, n5895, n5892, n5889, n5886, n5883, n5880, n5877, n5874, n5871, n5868, n5865, n5862, n5859, n5856, n5853, n5850, n5847, n5844, n5841, n5838, n5835, n5832, n5829, n5826, n5823, n5820, n5817, n5814, n5811, n5808, n5805, n5802, n5799, n5796, n5793, n5790, n5787, n5784, n5781, n5778, n5775, n5772, n5769, n5766, n5763, n5760, n5757, n5754, n5751, n5748, n5745, n5742, n5739, n5736, n5733, n5730, n5727, n5724, n5721, n5718, n5715, n5712, n5709, n5706, n5703, n5700, n5697, n5694, n5691, n5688, n5685, n5682, n5679, n5676, n5673, n5670, n5667, n5664, n5661, n5658, n5655, n5652, n5649, n5646, n5643, n5640, n5637, n5634, n5631, n5628, n5625, n5622, n5619, n5616, n5613, n5610, n5607, n5604, n5601, n5598, n5595, n5592, n5589, n5586, n5583, n5580, n5577, n5574, n5571, n5568, n5565, n5562, n5559, n5556, n5553, n5550, n5547, n5544, n5541, n5538, n5535, n5532, n5529, n5526, n5523, n5520, n5517, n5514, n5511, n5508, n5505, n5502, n5499, n5496, n5493, n5490, n5487, n5484, n5481, n5478, n5475, n5472, n5469, n5466, n5463, n5460, n5457, n5454, n5451, n5448, n5445, n5442, n5439, n5436, n5433, n5430, n5427, n5424, n5421, n5418, n5415, n5412, n5409, n5406, n5403, n5400, n5397, n5394, n5391, n5388, n5385, n5382, n5379, n5376, n5373, n5370, n5367, n5364, n5361, n5358, n5355, n5352, n5349, n5346, n5343, n5340, n5337, n5334, n5331, n5328, n5325, n5322, n5319, n5316, n5313, n5310, n5307, n5304, n5301, n5298, n5295, n5292, n5289, n5286, n5283, n5280, n5277, n5274, n5271, n5268, n5265, n5262, n5259, n5256, n5253, n5250, n5247, n5244, n5241, n5238, n5235, n5232, n5229, n5226, n5223, n5220, n5217, n5214, n5211, n5208, n5205, n5202, n5199, n5196, n5193, n5190, n5187, n5184, n5181, n5178, n5175, n5172, n5169, n5166, n5163, n5160, n5157, n5154, n5151, n5148, n5145, n5142, n5139, n5136, n5133, n5130, n5127, n5124, n5121, n5118, n5115, n5112, n5109, n5106, n5103, n5100, n5097, n5094, n5091, n5088, n5085, n5082, n5079, n5076, n5073, n5070, n5067, n5064, n5061, n5058, n5055, n5052, n5049, n5046, n5043, n5040, n5037, n5034, n5031, n5028, n5025, n5022, n5019, n5016, n5013, n5010, n5007, n5004, n5001, n4998, n4995, n4992, n4989, n4986, n4983, n4980, n4977, n4974, n4971, n4968, n4965, n4962, n4959, n4956, n4953, n4950, n4947, n4944, n4941, n4938, n4935, n4932, n4929, n4926, n4923, n4920, n4917, n4914, n4911, n4908, n4905, n4902, n4899, n4896, n4893, n4890, n4887, n4884, n4881, n4878, n4875, n4872, n4869, n4866, n4863, n4860, n4857, n4854, n4851, n4848, n4845, n4842, n4839, n4836, n4833, n4830, n4827, n4824, n4821, n4818, n4815, n4812, n4809, n4806, n4803, n4800, n4797, n4794, n4791, n4788, n4785, n4782, n4779, n4776, n4773, n4770, n4767, n4764, n4761, n4758, n4755, n4752, n4749, n4746, n4743, n4740, n4737, n4734, n4731, n4728, n4725, n4722, n4719, n4716, n4713, n4710, n4707, n4704, n4701, n4698, n4695, n4692, n4689, n4686, n4683, n4680, n4677, n4674, n4671, n4668, n4665, n4662, n4659, n4656, n4653, n4650, n4647, n4644, n4641, n4638, n4635, n4632, n4629, n4626, n4623, n4620, n4617, n4614, n4611, n4608, n4605, n4602, n4599, n4596, n4593, n4590, n4587, n4584, n4581, n4578, n4575, n4572, n4569, n4566, n4563, n4560, n4557, n4554, n4551, n4548, n4545, n4542, n4539, n4536, n4533, n4530, n4527, n4524, n4521, n4518, n4515, n4512, n4509, n4506, n4503, n4500, n4497, n4494, n4491, n4488, n4485, n4482, n4479, n4476, n4473, n4470, n4467, n4464, n4461, n4458, n4455, n4452, n4449, n4446, n4443, n4440, n4437, n4434, n4431, n4428, n4425, n4422, n4419, n4416, n4413, n4410, n4407, n4404, n4401, n4398, n4395, n4392, n4389, n4386, n4383, n4380, n4377, n4374, n4371, n4368, n4365};
  /* fppowtf32.vhdl:1117:4  */
  always @*
    case (n7436)
      1024'b1000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01111111111000;
      1024'b0100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01111111110000;
      1024'b0010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01111111101000;
      1024'b0001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01111111100000;
      1024'b0000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01111111011000;
      1024'b0000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01111111010000;
      1024'b0000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01111111001000;
      1024'b0000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01111111000000;
      1024'b0000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01111110111000;
      1024'b0000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01111110110000;
      1024'b0000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01111110101000;
      1024'b0000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01111110100001;
      1024'b0000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01111110011001;
      1024'b0000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01111110010001;
      1024'b0000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01111110001001;
      1024'b0000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01111110000001;
      1024'b0000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01111101111001;
      1024'b0000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01111101110001;
      1024'b0000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01111101101001;
      1024'b0000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01111101100010;
      1024'b0000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01111101011010;
      1024'b0000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01111101010010;
      1024'b0000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01111101001010;
      1024'b0000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01111101000010;
      1024'b0000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01111100111010;
      1024'b0000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01111100110011;
      1024'b0000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01111100101011;
      1024'b0000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01111100100011;
      1024'b0000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01111100011011;
      1024'b0000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01111100010011;
      1024'b0000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01111100001100;
      1024'b0000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01111100000100;
      1024'b0000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01111011111100;
      1024'b0000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01111011110100;
      1024'b0000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01111011101101;
      1024'b0000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01111011100101;
      1024'b0000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01111011011101;
      1024'b0000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01111011010110;
      1024'b0000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01111011001110;
      1024'b0000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01111011000110;
      1024'b0000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01111010111110;
      1024'b0000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01111010110111;
      1024'b0000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01111010101111;
      1024'b0000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01111010100111;
      1024'b0000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01111010100000;
      1024'b0000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01111010011000;
      1024'b0000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01111010010000;
      1024'b0000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01111010001001;
      1024'b0000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01111010000001;
      1024'b0000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01111001111010;
      1024'b0000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01111001110010;
      1024'b0000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01111001101010;
      1024'b0000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01111001100011;
      1024'b0000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01111001011011;
      1024'b0000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01111001010100;
      1024'b0000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01111001001100;
      1024'b0000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01111001000100;
      1024'b0000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01111000111101;
      1024'b0000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01111000110101;
      1024'b0000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01111000101110;
      1024'b0000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01111000100110;
      1024'b0000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01111000011111;
      1024'b0000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01111000010111;
      1024'b0000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01111000010000;
      1024'b0000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01111000001000;
      1024'b0000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01111000000001;
      1024'b0000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01110111111001;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01110111110010;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01110111101010;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01110111100011;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01110111011011;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01110111010100;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01110111001100;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01110111000101;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01110110111101;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01110110110110;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01110110101111;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01110110100111;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01110110100000;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01110110011000;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01110110010001;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01110110001010;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01110110000010;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01110101111011;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01110101110011;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01110101101100;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01110101100101;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01110101011101;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01110101010110;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01110101001111;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01110101000111;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01110101000000;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01110100111001;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01110100110001;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01110100101010;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01110100100011;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01110100011100;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01110100010100;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01110100001101;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01110100000110;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01110011111111;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01110011110111;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01110011110000;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01110011101001;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01110011100010;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01110011011010;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01110011010011;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01110011001100;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01110011000101;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01110010111110;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01110010110110;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01110010101111;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01110010101000;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01110010100001;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01110010011010;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01110010010011;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01110010001011;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01110010000100;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01110001111101;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01110001110110;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01110001101111;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01110001101000;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01110001100001;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01110001011010;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01110001010011;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01110001001100;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01110001000100;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01110000111101;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01110000110110;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01110000101111;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01110000101000;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01110000100001;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01110000011010;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01110000010011;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01110000001100;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01110000000101;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01101111111110;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01101111110111;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01101111110000;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01101111101001;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01101111100010;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01101111011011;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01101111010100;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01101111001101;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01101111000110;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01101110111111;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01101110111001;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01101110110010;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01101110101011;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01101110100100;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01101110011101;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01101110010110;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01101110001111;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01101110001000;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01101110000001;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01101101111010;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01101101110100;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01101101101101;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01101101100110;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01101101011111;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01101101011000;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01101101010001;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01101101001010;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01101101000100;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01101100111101;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01101100110110;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01101100101111;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01101100101000;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01101100100010;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01101100011011;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01101100010100;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01101100001101;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01101100000111;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01101100000000;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01101011111001;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01101011110010;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01101011101100;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01101011100101;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01101011011110;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01101011010111;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01101011010001;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01101011001010;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01101011000011;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01101010111101;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01101010110110;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01101010101111;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01101010101001;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01101010100010;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01101010011011;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01101010010101;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01101010001110;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01101010000111;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01101010000001;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01101001111010;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01101001110100;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01101001101101;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01101001100110;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01101001100000;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01101001011001;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01101001010011;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01101001001100;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01101001000101;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01101000111111;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01101000111000;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01101000110010;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01101000101011;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01101000100101;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01101000011110;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01101000011000;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01101000010001;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01101000001011;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01101000000100;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01100111111110;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01100111110111;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01100111110001;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01100111101010;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01100111100100;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01100111011101;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01100111010111;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01100111010000;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01100111001010;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01100111000011;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01100110111101;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01100110110110;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01100110110000;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01100110101010;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01100110100011;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01100110011101;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01100110010110;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01100110010000;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01100110001010;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01100110000011;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01100101111101;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01100101110110;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01100101110000;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01100101101010;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01100101100011;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01100101011101;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01100101010111;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01100101010000;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01100101001010;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01100101000100;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01100100111101;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01100100110111;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01100100110001;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01100100101011;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01100100100100;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01100100011110;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01100100011000;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01100100010001;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01100100001011;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01100100000101;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01100011111111;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01100011111000;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01100011110010;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01100011101100;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01100011100110;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01100011011111;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01100011011001;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01100011010011;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01100011001101;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01100011000111;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01100011000000;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01100010111010;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01100010110100;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01100010101110;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01100010101000;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01100010100010;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01100010011011;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01100010010101;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01100010001111;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01100010001001;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01100010000011;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01100001111101;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01100001110111;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01100001110001;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01100001101010;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01100001100100;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01100001011110;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01100001011000;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01100001010010;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01100001001100;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01100001000110;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01100001000000;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01100000111010;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01100000110100;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01100000101110;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01100000101000;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01100000100010;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01100000011100;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01100000010110;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01100000010000;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01100000001010;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01100000000100;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01011111111110;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01011111111000;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01011111110010;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01011111101100;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01011111100110;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01011111100000;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01011111011010;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01011111010100;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01011111001110;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01011111001000;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01011111000010;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01011110111100;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01011110110110;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01011110110000;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01011110101010;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01011110100100;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01011110011110;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01011110011000;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01011110010011;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01011110001101;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01011110000111;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01011110000001;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01011101111011;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01011101110101;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01011101101111;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01011101101001;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01011101100100;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01011101011110;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01011101011000;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01011101010010;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01011101001100;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01011101000110;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01011101000001;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01011100111011;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01011100110101;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01011100101111;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01011100101001;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01011100100100;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01011100011110;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01011100011000;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01011100010010;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01011100001100;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01011100000111;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01011100000001;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01011011111011;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01011011110101;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01011011110000;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01011011101010;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01011011100100;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01011011011111;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01011011011001;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01011011010011;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01011011001101;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01011011001000;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01011011000010;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01011010111100;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01011010110111;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01011010110001;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01011010101011;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01011010100110;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01011010100000;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01011010011010;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01011010010101;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01011010001111;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01011010001001;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01011010000100;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01011001111110;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01011001111001;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01011001110011;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01011001101101;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01011001101000;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01011001100010;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01011001011101;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01011001010111;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01011001010001;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01011001001100;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01011001000110;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01011001000001;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01011000111011;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01011000110110;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01011000110000;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01011000101010;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01011000100101;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01011000011111;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01011000011010;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01011000010100;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01011000001111;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01011000001001;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01011000000100;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01010111111110;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01010111111001;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01010111110011;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01010111101110;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01010111101000;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01010111100011;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01010111011101;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01010111011000;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01010111010010;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01010111001101;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01010111001000;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01010111000010;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01010110111101;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01010110110111;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01010110110010;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01010110101100;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01010110100111;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01010110100010;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01010110011100;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01010110010111;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01010110010001;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01010110001100;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01010110000111;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01010110000001;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01010101111100;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01010101110110;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01010101110001;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01010101101100;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01010101100110;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01010101100001;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01010101011100;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01010101010110;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01010101010001;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01010101001100;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01010101000110;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01010101000001;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01010100111100;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01010100110110;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01010100110001;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01010100101100;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01010100100111;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01010100100001;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01010100011100;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01010100010111;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01010100010001;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01010100001100;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01010100000111;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01010100000010;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01010011111100;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01010011110111;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01010011110010;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01010011101101;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01010011100111;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01010011100010;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01010011011101;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01010011011000;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01010011010011;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01010011001101;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01010011001000;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01010011000011;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01010010111110;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01010010111001;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01010010110011;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01010010101110;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01010010101001;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01010010100100;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01010010011111;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01010010011010;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01010010010101;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01010010001111;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01010010001010;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01010010000101;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01010010000000;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01010001111011;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01010001110110;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01010001110001;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01010001101100;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01010001100110;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01010001100001;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01010001011100;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01010001010111;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01010001010010;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01010001001101;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01010001001000;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01010001000011;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01010000111110;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01010000111001;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01010000110100;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01010000101111;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01010000101010;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01010000100101;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01010000100000;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01010000011010;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01010000010101;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01010000010000;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01010000001011;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01010000000110;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01010000000001;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01001111111100;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01001111110111;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01001111110010;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01001111101101;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01001111101000;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01001111100011;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01001111011111;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01001111011010;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01001111010101;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01001111010000;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01001111001011;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01001111000110;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01001111000001;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01001110111100;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01001110110111;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01001110110010;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01001110101101;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01001110101000;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01001110100011;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01001110011110;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01001110011001;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01001110010101;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01001110010000;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01001110001011;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01001110000110;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01001110000001;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01001101111100;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01001101110111;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01001101110010;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01001101101110;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b01001101101001;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b11010010110101;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b11010010101000;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b11010010011011;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b11010010001110;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b11010010000001;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b11010001110011;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b11010001100110;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b11010001011001;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b11010001001100;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b11010000111111;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b11010000110010;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b11010000100101;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b11010000011000;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b11010000001011;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b11001111111110;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b11001111110001;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b11001111100100;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b11001111010111;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b11001111001010;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b11001110111101;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b11001110110000;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b11001110100011;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b11001110010110;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b11001110001001;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b11001101111101;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b11001101110000;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b11001101100011;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b11001101010110;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b11001101001001;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b11001100111100;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b11001100110000;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b11001100100011;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b11001100010110;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b11001100001001;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b11001011111100;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b11001011110000;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b11001011100011;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b11001011010110;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b11001011001010;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b11001010111101;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b11001010110000;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b11001010100100;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b11001010010111;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b11001010001010;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b11001001111110;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b11001001110001;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b11001001100100;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b11001001011000;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b11001001001011;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b11001000111111;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b11001000110010;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b11001000100110;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b11001000011001;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b11001000001101;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b11001000000000;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b11000111110100;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b11000111100111;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b11000111011011;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b11000111001110;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b11000111000010;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b11000110110101;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b11000110101001;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b11000110011100;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b11000110010000;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b11000110000100;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b11000101110111;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b11000101101011;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b11000101011111;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b11000101010010;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b11000101000110;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b11000100111010;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b11000100101101;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b11000100100001;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b11000100010101;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b11000100001000;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b11000011111100;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b11000011110000;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b11000011100100;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b11000011011000;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b11000011001011;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b11000010111111;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b11000010110011;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b11000010100111;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b11000010011011;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b11000010001110;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b11000010000010;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b11000001110110;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b11000001101010;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b11000001011110;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b11000001010010;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b11000001000110;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b11000000111010;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b11000000101110;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b11000000100010;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b11000000010110;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b11000000001010;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b10111111111110;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b10111111110010;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b10111111100110;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b10111111011010;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b10111111001110;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b10111111000010;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b10111110110110;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b10111110101010;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b10111110011110;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b10111110010010;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b10111110000110;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b10111101111010;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b10111101101111;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b10111101100011;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b10111101010111;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b10111101001011;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b10111100111111;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b10111100110011;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b10111100101000;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b10111100011100;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b10111100010000;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b10111100000100;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b10111011111001;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b10111011101101;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b10111011100001;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b10111011010101;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b10111011001010;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b10111010111110;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b10111010110010;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b10111010100111;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b10111010011011;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b10111010001111;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b10111010000100;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b10111001111000;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b10111001101100;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b10111001100001;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b10111001010101;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b10111001001010;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b10111000111110;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b10111000110011;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b10111000100111;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b10111000011011;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b10111000010000;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b10111000000100;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b10110111111001;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b10110111101101;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b10110111100010;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b10110111010110;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b10110111001011;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b10110111000000;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b10110110110100;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b10110110101001;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b10110110011101;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b10110110010010;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b10110110000111;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b10110101111011;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b10110101110000;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b10110101100100;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b10110101011001;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b10110101001110;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b10110101000010;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b10110100110111;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b10110100101100;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b10110100100001;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b10110100010101;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b10110100001010;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b10110011111111;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b10110011110100;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b10110011101000;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b10110011011101;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b10110011010010;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b10110011000111;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b10110010111011;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b10110010110000;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b10110010100101;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b10110010011010;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b10110010001111;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b10110010000100;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b10110001111001;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b10110001101101;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b10110001100010;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b10110001010111;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b10110001001100;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b10110001000001;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b10110000110110;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b10110000101011;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b10110000100000;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b10110000010101;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b10110000001010;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b10101111111111;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b10101111110100;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b10101111101001;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b10101111011110;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b10101111010011;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b10101111001000;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b10101110111101;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b10101110110010;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b10101110100111;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b10101110011100;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b10101110010001;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b10101110000111;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b10101101111100;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b10101101110001;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b10101101100110;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b10101101011011;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b10101101010000;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b10101101000101;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b10101100111011;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b10101100110000;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b10101100100101;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b10101100011010;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b10101100010000;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b10101100000101;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b10101011111010;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b10101011101111;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b10101011100101;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b10101011011010;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b10101011001111;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b10101011000100;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b10101010111010;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b10101010101111;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b10101010100100;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b10101010011010;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b10101010001111;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b10101010000100;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b10101001111010;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b10101001101111;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b10101001100101;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b10101001011010;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b10101001001111;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b10101001000101;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b10101000111010;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b10101000110000;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b10101000100101;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b10101000011011;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b10101000010000;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b10101000000110;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b10100111111011;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b10100111110001;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b10100111100110;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b10100111011100;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b10100111010001;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b10100111000111;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b10100110111100;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b10100110110010;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b10100110101000;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b10100110011101;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b10100110010011;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b10100110001000;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b10100101111110;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b10100101110100;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b10100101101001;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b10100101011111;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b10100101010101;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b10100101001010;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b10100101000000;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b10100100110110;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b10100100101011;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b10100100100001;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b10100100010111;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b10100100001100;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b10100100000010;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b10100011111000;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b10100011101110;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b10100011100100;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b10100011011001;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b10100011001111;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b10100011000101;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b10100010111011;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b10100010110001;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b10100010100110;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b10100010011100;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b10100010010010;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b10100010001000;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b10100001111110;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b10100001110100;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b10100001101010;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b10100001011111;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b10100001010101;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b10100001001011;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b10100001000001;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b10100000110111;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b10100000101101;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b10100000100011;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b10100000011001;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b10100000001111;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b10100000000101;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b10011111111011;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b10011111110001;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b10011111100111;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b10011111011101;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b10011111010011;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b10011111001001;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b10011110111111;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b10011110110101;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b10011110101011;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b10011110100001;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b10011110011000;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b10011110001110;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b10011110000100;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b10011101111010;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b10011101110000;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b10011101100110;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b10011101011100;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b10011101010010;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b10011101001001;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b10011100111111;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b10011100110101;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b10011100101011;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b10011100100001;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b10011100011000;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b10011100001110;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b10011100000100;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b10011011111010;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b10011011110001;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b10011011100111;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b10011011011101;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b10011011010100;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b10011011001010;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b10011011000000;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b10011010110110;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b10011010101101;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b10011010100011;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b10011010011001;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b10011010010000;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b10011010000110;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b10011001111101;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b10011001110011;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b10011001101001;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b10011001100000;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b10011001010110;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b10011001001101;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b10011001000011;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b10011000111001;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b10011000110000;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b10011000100110;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b10011000011101;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b10011000010011;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b10011000001010;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b10011000000000;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b10010111110111;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b10010111101101;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b10010111100100;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b10010111011010;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b10010111010001;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b10010111000111;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b10010110111110;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b10010110110101;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b10010110101011;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b10010110100010;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b10010110011000;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b10010110001111;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b10010110000110;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b10010101111100;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b10010101110011;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b10010101101001;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b10010101100000;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b10010101010111;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b10010101001101;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b10010101000100;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b10010100111011;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b10010100110001;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b10010100101000;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b10010100011111;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b10010100010110;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b10010100001100;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b10010100000011;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b10010011111010;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b10010011110001;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b10010011100111;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b10010011011110;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b10010011010101;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b10010011001100;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b10010011000011;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b10010010111001;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b10010010110000;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b10010010100111;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b10010010011110;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b10010010010101;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b10010010001100;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b10010010000010;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b10010001111001;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b10010001110000;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b10010001100111;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b10010001011110;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b10010001010101;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b10010001001100;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b10010001000011;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b10010000111010;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b10010000110001;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b10010000101000;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b10010000011111;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b10010000010110;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b10010000001101;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b10010000000100;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b10001111111011;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b10001111110010;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b10001111101001;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b10001111100000;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b10001111010111;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b10001111001110;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b10001111000101;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b10001110111100;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b10001110110011;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b10001110101010;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b10001110100001;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b10001110011000;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b10001110001111;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b10001110000110;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b10001101111101;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b10001101110101;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b10001101101100;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b10001101100011;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b10001101011010;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b10001101010001;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b10001101001000;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b10001101000000;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b10001100110111;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b10001100101110;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b10001100100101;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b10001100011100;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b10001100010100;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b10001100001011;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b10001100000010;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b10001011111001;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b10001011110001;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b10001011101000;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b10001011011111;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b10001011010110;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b10001011001110;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b10001011000101;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b10001010111100;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b10001010110100;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b10001010101011;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b10001010100010;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b10001010011010;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b10001010010001;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b10001010001000;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b10001010000000;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b10001001110111;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b10001001101111;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b10001001100110;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b10001001011101;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b10001001010101;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b10001001001100;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b10001001000100;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b10001000111011;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b10001000110010;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b10001000101010;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b10001000100001;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b10001000011001;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b10001000010000;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b10001000001000;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b10000111111111;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b10000111110111;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000: n7437 = 14'b10000111101110;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000: n7437 = 14'b10000111100110;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000: n7437 = 14'b10000111011101;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000: n7437 = 14'b10000111010101;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000: n7437 = 14'b10000111001100;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000: n7437 = 14'b10000111000100;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000: n7437 = 14'b10000110111100;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000: n7437 = 14'b10000110110011;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000: n7437 = 14'b10000110101011;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000: n7437 = 14'b10000110100010;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000: n7437 = 14'b10000110011010;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000: n7437 = 14'b10000110010010;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000: n7437 = 14'b10000110001001;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000: n7437 = 14'b10000110000001;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000: n7437 = 14'b10000101111000;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000: n7437 = 14'b10000101110000;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000: n7437 = 14'b10000101101000;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000: n7437 = 14'b10000101011111;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000: n7437 = 14'b10000101010111;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000: n7437 = 14'b10000101001111;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000: n7437 = 14'b10000101000110;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000: n7437 = 14'b10000100111110;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000: n7437 = 14'b10000100110110;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000: n7437 = 14'b10000100101101;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000: n7437 = 14'b10000100100101;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000: n7437 = 14'b10000100011101;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000: n7437 = 14'b10000100010101;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000: n7437 = 14'b10000100001100;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000: n7437 = 14'b10000100000100;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000: n7437 = 14'b10000011111100;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000: n7437 = 14'b10000011110100;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000: n7437 = 14'b10000011101011;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000: n7437 = 14'b10000011100011;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000: n7437 = 14'b10000011011011;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000: n7437 = 14'b10000011010011;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000: n7437 = 14'b10000011001010;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000: n7437 = 14'b10000011000010;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000: n7437 = 14'b10000010111010;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000: n7437 = 14'b10000010110010;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000: n7437 = 14'b10000010101010;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000: n7437 = 14'b10000010100010;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000: n7437 = 14'b10000010011001;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000: n7437 = 14'b10000010010001;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000: n7437 = 14'b10000010001001;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000: n7437 = 14'b10000010000001;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000: n7437 = 14'b10000001111001;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000: n7437 = 14'b10000001110001;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000: n7437 = 14'b10000001101001;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000: n7437 = 14'b10000001100001;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000: n7437 = 14'b10000001011000;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000: n7437 = 14'b10000001010000;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000: n7437 = 14'b10000001001000;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000: n7437 = 14'b10000001000000;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000: n7437 = 14'b10000000111000;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000: n7437 = 14'b10000000110000;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000: n7437 = 14'b10000000101000;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000: n7437 = 14'b10000000100000;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000: n7437 = 14'b10000000011000;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100: n7437 = 14'b10000000010000;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010: n7437 = 14'b10000000001000;
      1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001: n7437 = 14'b10000000000000;
      default: n7437 = 14'bX;
    endcase
endmodule

module intadder_13_freq500_uid102
  (input  clk,
   input  [12:0] x,
   input  [12:0] y,
   input  cin,
   output [12:0] r);
  wire [12:0] rtmp;
  wire [12:0] x_d1;
  wire [12:0] x_d2;
  wire [12:0] x_d3;
  wire [12:0] y_d1;
  wire cin_d1;
  wire cin_d2;
  wire cin_d3;
  wire cin_d4;
  wire cin_d5;
  wire cin_d6;
  wire cin_d7;
  wire cin_d8;
  wire cin_d9;
  wire cin_d10;
  wire cin_d11;
  wire cin_d12;
  wire cin_d13;
  wire cin_d14;
  wire cin_d15;
  wire cin_d16;
  wire cin_d17;
  wire cin_d18;
  wire [12:0] n4337;
  wire [12:0] n4338;
  wire [12:0] n4339;
  reg [12:0] n4340;
  reg [12:0] n4341;
  reg [12:0] n4342;
  reg [12:0] n4343;
  reg n4344;
  reg n4345;
  reg n4346;
  reg n4347;
  reg n4348;
  reg n4349;
  reg n4350;
  reg n4351;
  reg n4352;
  reg n4353;
  reg n4354;
  reg n4355;
  reg n4356;
  reg n4357;
  reg n4358;
  reg n4359;
  reg n4360;
  reg n4361;
  assign r = rtmp; //(module output)
  /* fppowtf32.vhdl:4953:8  */
  assign rtmp = n4339; // (signal)
  /* fppowtf32.vhdl:4955:8  */
  assign x_d1 = n4340; // (signal)
  /* fppowtf32.vhdl:4955:14  */
  assign x_d2 = n4341; // (signal)
  /* fppowtf32.vhdl:4955:20  */
  assign x_d3 = n4342; // (signal)
  /* fppowtf32.vhdl:4957:8  */
  assign y_d1 = n4343; // (signal)
  /* fppowtf32.vhdl:4959:8  */
  assign cin_d1 = n4344; // (signal)
  /* fppowtf32.vhdl:4959:16  */
  assign cin_d2 = n4345; // (signal)
  /* fppowtf32.vhdl:4959:24  */
  assign cin_d3 = n4346; // (signal)
  /* fppowtf32.vhdl:4959:32  */
  assign cin_d4 = n4347; // (signal)
  /* fppowtf32.vhdl:4959:40  */
  assign cin_d5 = n4348; // (signal)
  /* fppowtf32.vhdl:4959:48  */
  assign cin_d6 = n4349; // (signal)
  /* fppowtf32.vhdl:4959:56  */
  assign cin_d7 = n4350; // (signal)
  /* fppowtf32.vhdl:4959:64  */
  assign cin_d8 = n4351; // (signal)
  /* fppowtf32.vhdl:4959:72  */
  assign cin_d9 = n4352; // (signal)
  /* fppowtf32.vhdl:4959:80  */
  assign cin_d10 = n4353; // (signal)
  /* fppowtf32.vhdl:4959:89  */
  assign cin_d11 = n4354; // (signal)
  /* fppowtf32.vhdl:4959:98  */
  assign cin_d12 = n4355; // (signal)
  /* fppowtf32.vhdl:4959:107  */
  assign cin_d13 = n4356; // (signal)
  /* fppowtf32.vhdl:4959:116  */
  assign cin_d14 = n4357; // (signal)
  /* fppowtf32.vhdl:4959:125  */
  assign cin_d15 = n4358; // (signal)
  /* fppowtf32.vhdl:4959:134  */
  assign cin_d16 = n4359; // (signal)
  /* fppowtf32.vhdl:4959:143  */
  assign cin_d17 = n4360; // (signal)
  /* fppowtf32.vhdl:4959:152  */
  assign cin_d18 = n4361; // (signal)
  /* fppowtf32.vhdl:4989:17  */
  assign n4337 = x_d3 + y_d1;
  /* fppowtf32.vhdl:4989:24  */
  assign n4338 = {12'b0, cin_d18};  //  uext
  /* fppowtf32.vhdl:4989:24  */
  assign n4339 = n4337 + n4338;
  /* fppowtf32.vhdl:4964:10  */
  always @(posedge clk)
    n4340 <= x;
  /* fppowtf32.vhdl:4964:10  */
  always @(posedge clk)
    n4341 <= x_d1;
  /* fppowtf32.vhdl:4964:10  */
  always @(posedge clk)
    n4342 <= x_d2;
  /* fppowtf32.vhdl:4964:10  */
  always @(posedge clk)
    n4343 <= y;
  /* fppowtf32.vhdl:4964:10  */
  always @(posedge clk)
    n4344 <= cin;
  /* fppowtf32.vhdl:4964:10  */
  always @(posedge clk)
    n4345 <= cin_d1;
  /* fppowtf32.vhdl:4964:10  */
  always @(posedge clk)
    n4346 <= cin_d2;
  /* fppowtf32.vhdl:4964:10  */
  always @(posedge clk)
    n4347 <= cin_d3;
  /* fppowtf32.vhdl:4964:10  */
  always @(posedge clk)
    n4348 <= cin_d4;
  /* fppowtf32.vhdl:4964:10  */
  always @(posedge clk)
    n4349 <= cin_d5;
  /* fppowtf32.vhdl:4964:10  */
  always @(posedge clk)
    n4350 <= cin_d6;
  /* fppowtf32.vhdl:4964:10  */
  always @(posedge clk)
    n4351 <= cin_d7;
  /* fppowtf32.vhdl:4964:10  */
  always @(posedge clk)
    n4352 <= cin_d8;
  /* fppowtf32.vhdl:4964:10  */
  always @(posedge clk)
    n4353 <= cin_d9;
  /* fppowtf32.vhdl:4964:10  */
  always @(posedge clk)
    n4354 <= cin_d10;
  /* fppowtf32.vhdl:4964:10  */
  always @(posedge clk)
    n4355 <= cin_d11;
  /* fppowtf32.vhdl:4964:10  */
  always @(posedge clk)
    n4356 <= cin_d12;
  /* fppowtf32.vhdl:4964:10  */
  always @(posedge clk)
    n4357 <= cin_d13;
  /* fppowtf32.vhdl:4964:10  */
  always @(posedge clk)
    n4358 <= cin_d14;
  /* fppowtf32.vhdl:4964:10  */
  always @(posedge clk)
    n4359 <= cin_d15;
  /* fppowtf32.vhdl:4964:10  */
  always @(posedge clk)
    n4360 <= cin_d16;
  /* fppowtf32.vhdl:4964:10  */
  always @(posedge clk)
    n4361 <= cin_d17;
endmodule

module fixrealkcm_freq500_uid89
  (input  clk,
   input  [7:0] x,
   output [20:0] r);
  wire [4:0] fixrealkcm_freq500_uid89_a0;
  wire [20:0] fixrealkcm_freq500_uid89_t0;
  wire [20:0] fixrealkcm_freq500_uid89_t0_copy93;
  wire bh90_w0_0;
  wire bh90_w1_0;
  wire bh90_w2_0;
  wire bh90_w3_0;
  wire bh90_w4_0;
  wire bh90_w5_0;
  wire bh90_w6_0;
  wire bh90_w7_0;
  wire bh90_w8_0;
  wire bh90_w9_0;
  wire bh90_w10_0;
  wire bh90_w11_0;
  wire bh90_w12_0;
  wire bh90_w13_0;
  wire bh90_w14_0;
  wire bh90_w15_0;
  wire bh90_w16_0;
  wire bh90_w17_0;
  wire bh90_w18_0;
  wire bh90_w19_0;
  wire bh90_w20_0;
  wire [2:0] fixrealkcm_freq500_uid89_a1;
  wire [15:0] fixrealkcm_freq500_uid89_t1;
  wire [15:0] fixrealkcm_freq500_uid89_t1_copy96;
  wire bh90_w0_1;
  wire bh90_w1_1;
  wire bh90_w2_1;
  wire bh90_w3_1;
  wire bh90_w4_1;
  wire bh90_w5_1;
  wire bh90_w6_1;
  wire bh90_w7_1;
  wire bh90_w8_1;
  wire bh90_w9_1;
  wire bh90_w10_1;
  wire bh90_w11_1;
  wire bh90_w12_1;
  wire bh90_w13_1;
  wire bh90_w14_1;
  wire bh90_w15_1;
  wire [20:0] bitheapfinaladd_bh90_in0;
  wire [20:0] bitheapfinaladd_bh90_in1;
  wire bitheapfinaladd_bh90_cin;
  wire [20:0] bitheapfinaladd_bh90_out;
  wire [20:0] bitheapresult_bh90;
  wire [20:0] outres;
  wire [4:0] n4223;
  wire [20:0] fixrealkcm_freq500_uid89_table0_n4224;
  wire n4227;
  wire n4228;
  wire n4229;
  wire n4230;
  wire n4231;
  wire n4232;
  wire n4233;
  wire n4234;
  wire n4235;
  wire n4236;
  wire n4237;
  wire n4238;
  wire n4239;
  wire n4240;
  wire n4241;
  wire n4242;
  wire n4243;
  wire n4244;
  wire n4245;
  wire n4246;
  wire n4247;
  wire [2:0] n4248;
  wire [15:0] fixrealkcm_freq500_uid89_table1_n4249;
  wire n4252;
  wire n4253;
  wire n4254;
  wire n4255;
  wire n4256;
  wire n4257;
  wire n4258;
  wire n4259;
  wire n4260;
  wire n4261;
  wire n4262;
  wire n4263;
  wire n4264;
  wire n4265;
  wire n4266;
  wire n4267;
  wire [1:0] n4269;
  wire [2:0] n4270;
  wire [3:0] n4271;
  wire [4:0] n4272;
  wire [5:0] n4273;
  wire [6:0] n4274;
  wire [7:0] n4275;
  wire [8:0] n4276;
  wire [9:0] n4277;
  wire [10:0] n4278;
  wire [11:0] n4279;
  wire [12:0] n4280;
  wire [13:0] n4281;
  wire [14:0] n4282;
  wire [15:0] n4283;
  wire [16:0] n4284;
  wire [17:0] n4285;
  wire [18:0] n4286;
  wire [19:0] n4287;
  wire [20:0] n4288;
  wire [5:0] n4290;
  wire [6:0] n4291;
  wire [7:0] n4292;
  wire [8:0] n4293;
  wire [9:0] n4294;
  wire [10:0] n4295;
  wire [11:0] n4296;
  wire [12:0] n4297;
  wire [13:0] n4298;
  wire [14:0] n4299;
  wire [15:0] n4300;
  wire [16:0] n4301;
  wire [17:0] n4302;
  wire [18:0] n4303;
  wire [19:0] n4304;
  wire [20:0] n4305;
  wire [20:0] bitheapfinaladd_bh90_n4307;
  assign r = outres; //(module output)
  /* fppowtf32.vhdl:4754:8  */
  assign fixrealkcm_freq500_uid89_a0 = n4223; // (signal)
  /* fppowtf32.vhdl:4756:8  */
  assign fixrealkcm_freq500_uid89_t0 = fixrealkcm_freq500_uid89_t0_copy93; // (signal)
  /* fppowtf32.vhdl:4758:8  */
  assign fixrealkcm_freq500_uid89_t0_copy93 = fixrealkcm_freq500_uid89_table0_n4224; // (signal)
  /* fppowtf32.vhdl:4760:8  */
  assign bh90_w0_0 = n4227; // (signal)
  /* fppowtf32.vhdl:4762:8  */
  assign bh90_w1_0 = n4228; // (signal)
  /* fppowtf32.vhdl:4764:8  */
  assign bh90_w2_0 = n4229; // (signal)
  /* fppowtf32.vhdl:4766:8  */
  assign bh90_w3_0 = n4230; // (signal)
  /* fppowtf32.vhdl:4768:8  */
  assign bh90_w4_0 = n4231; // (signal)
  /* fppowtf32.vhdl:4770:8  */
  assign bh90_w5_0 = n4232; // (signal)
  /* fppowtf32.vhdl:4772:8  */
  assign bh90_w6_0 = n4233; // (signal)
  /* fppowtf32.vhdl:4774:8  */
  assign bh90_w7_0 = n4234; // (signal)
  /* fppowtf32.vhdl:4776:8  */
  assign bh90_w8_0 = n4235; // (signal)
  /* fppowtf32.vhdl:4778:8  */
  assign bh90_w9_0 = n4236; // (signal)
  /* fppowtf32.vhdl:4780:8  */
  assign bh90_w10_0 = n4237; // (signal)
  /* fppowtf32.vhdl:4782:8  */
  assign bh90_w11_0 = n4238; // (signal)
  /* fppowtf32.vhdl:4784:8  */
  assign bh90_w12_0 = n4239; // (signal)
  /* fppowtf32.vhdl:4786:8  */
  assign bh90_w13_0 = n4240; // (signal)
  /* fppowtf32.vhdl:4788:8  */
  assign bh90_w14_0 = n4241; // (signal)
  /* fppowtf32.vhdl:4790:8  */
  assign bh90_w15_0 = n4242; // (signal)
  /* fppowtf32.vhdl:4792:8  */
  assign bh90_w16_0 = n4243; // (signal)
  /* fppowtf32.vhdl:4794:8  */
  assign bh90_w17_0 = n4244; // (signal)
  /* fppowtf32.vhdl:4796:8  */
  assign bh90_w18_0 = n4245; // (signal)
  /* fppowtf32.vhdl:4798:8  */
  assign bh90_w19_0 = n4246; // (signal)
  /* fppowtf32.vhdl:4906:35  */
  assign bh90_w20_0 = n4247; // (signal)
  /* fppowtf32.vhdl:4802:8  */
  assign fixrealkcm_freq500_uid89_a1 = n4248; // (signal)
  /* fppowtf32.vhdl:4804:8  */
  assign fixrealkcm_freq500_uid89_t1 = fixrealkcm_freq500_uid89_t1_copy96; // (signal)
  /* fppowtf32.vhdl:4806:8  */
  assign fixrealkcm_freq500_uid89_t1_copy96 = fixrealkcm_freq500_uid89_table1_n4249; // (signal)
  /* fppowtf32.vhdl:4808:8  */
  assign bh90_w0_1 = n4252; // (signal)
  /* fppowtf32.vhdl:4810:8  */
  assign bh90_w1_1 = n4253; // (signal)
  /* fppowtf32.vhdl:4812:8  */
  assign bh90_w2_1 = n4254; // (signal)
  /* fppowtf32.vhdl:4814:8  */
  assign bh90_w3_1 = n4255; // (signal)
  /* fppowtf32.vhdl:4816:8  */
  assign bh90_w4_1 = n4256; // (signal)
  /* fppowtf32.vhdl:4818:8  */
  assign bh90_w5_1 = n4257; // (signal)
  /* fppowtf32.vhdl:4820:8  */
  assign bh90_w6_1 = n4258; // (signal)
  /* fppowtf32.vhdl:4822:8  */
  assign bh90_w7_1 = n4259; // (signal)
  /* fppowtf32.vhdl:4824:8  */
  assign bh90_w8_1 = n4260; // (signal)
  /* fppowtf32.vhdl:4826:8  */
  assign bh90_w9_1 = n4261; // (signal)
  /* fppowtf32.vhdl:4828:8  */
  assign bh90_w10_1 = n4262; // (signal)
  /* fppowtf32.vhdl:4830:8  */
  assign bh90_w11_1 = n4263; // (signal)
  /* fppowtf32.vhdl:4832:8  */
  assign bh90_w12_1 = n4264; // (signal)
  /* fppowtf32.vhdl:4834:8  */
  assign bh90_w13_1 = n4265; // (signal)
  /* fppowtf32.vhdl:4836:8  */
  assign bh90_w14_1 = n4266; // (signal)
  /* fppowtf32.vhdl:4838:8  */
  assign bh90_w15_1 = n4267; // (signal)
  /* fppowtf32.vhdl:4840:8  */
  assign bitheapfinaladd_bh90_in0 = n4288; // (signal)
  /* fppowtf32.vhdl:4842:8  */
  assign bitheapfinaladd_bh90_in1 = n4305; // (signal)
  /* fppowtf32.vhdl:4844:8  */
  assign bitheapfinaladd_bh90_cin = 1'b0; // (signal)
  /* fppowtf32.vhdl:4846:8  */
  assign bitheapfinaladd_bh90_out = bitheapfinaladd_bh90_n4307; // (signal)
  /* fppowtf32.vhdl:4848:8  */
  assign bitheapresult_bh90 = bitheapfinaladd_bh90_out; // (signal)
  /* fppowtf32.vhdl:4850:8  */
  assign outres = bitheapresult_bh90; // (signal)
  /* fppowtf32.vhdl:4854:36  */
  assign n4223 = x[7:3]; // extract
  /* fppowtf32.vhdl:4855:4  */
  fixrealkcm_freq500_uid89_t0_freq500_uid92 fixrealkcm_freq500_uid89_table0 (
    .x(fixrealkcm_freq500_uid89_a0),
    .y(fixrealkcm_freq500_uid89_table0_n4224));
  /* fppowtf32.vhdl:4859:44  */
  assign n4227 = fixrealkcm_freq500_uid89_t0[0]; // extract
  /* fppowtf32.vhdl:4860:44  */
  assign n4228 = fixrealkcm_freq500_uid89_t0[1]; // extract
  /* fppowtf32.vhdl:4861:44  */
  assign n4229 = fixrealkcm_freq500_uid89_t0[2]; // extract
  /* fppowtf32.vhdl:4862:44  */
  assign n4230 = fixrealkcm_freq500_uid89_t0[3]; // extract
  /* fppowtf32.vhdl:4863:44  */
  assign n4231 = fixrealkcm_freq500_uid89_t0[4]; // extract
  /* fppowtf32.vhdl:4864:44  */
  assign n4232 = fixrealkcm_freq500_uid89_t0[5]; // extract
  /* fppowtf32.vhdl:4865:44  */
  assign n4233 = fixrealkcm_freq500_uid89_t0[6]; // extract
  /* fppowtf32.vhdl:4866:44  */
  assign n4234 = fixrealkcm_freq500_uid89_t0[7]; // extract
  /* fppowtf32.vhdl:4867:44  */
  assign n4235 = fixrealkcm_freq500_uid89_t0[8]; // extract
  /* fppowtf32.vhdl:4868:44  */
  assign n4236 = fixrealkcm_freq500_uid89_t0[9]; // extract
  /* fppowtf32.vhdl:4869:45  */
  assign n4237 = fixrealkcm_freq500_uid89_t0[10]; // extract
  /* fppowtf32.vhdl:4870:45  */
  assign n4238 = fixrealkcm_freq500_uid89_t0[11]; // extract
  /* fppowtf32.vhdl:4871:45  */
  assign n4239 = fixrealkcm_freq500_uid89_t0[12]; // extract
  /* fppowtf32.vhdl:4872:45  */
  assign n4240 = fixrealkcm_freq500_uid89_t0[13]; // extract
  /* fppowtf32.vhdl:4873:45  */
  assign n4241 = fixrealkcm_freq500_uid89_t0[14]; // extract
  /* fppowtf32.vhdl:4874:45  */
  assign n4242 = fixrealkcm_freq500_uid89_t0[15]; // extract
  /* fppowtf32.vhdl:4875:45  */
  assign n4243 = fixrealkcm_freq500_uid89_t0[16]; // extract
  /* fppowtf32.vhdl:4876:45  */
  assign n4244 = fixrealkcm_freq500_uid89_t0[17]; // extract
  /* fppowtf32.vhdl:4877:45  */
  assign n4245 = fixrealkcm_freq500_uid89_t0[18]; // extract
  /* fppowtf32.vhdl:4878:45  */
  assign n4246 = fixrealkcm_freq500_uid89_t0[19]; // extract
  /* fppowtf32.vhdl:4879:45  */
  assign n4247 = fixrealkcm_freq500_uid89_t0[20]; // extract
  /* fppowtf32.vhdl:4880:36  */
  assign n4248 = x[2:0]; // extract
  /* fppowtf32.vhdl:4881:4  */
  fixrealkcm_freq500_uid89_t1_freq500_uid95 fixrealkcm_freq500_uid89_table1 (
    .x(fixrealkcm_freq500_uid89_a1),
    .y(fixrealkcm_freq500_uid89_table1_n4249));
  /* fppowtf32.vhdl:4885:44  */
  assign n4252 = fixrealkcm_freq500_uid89_t1[0]; // extract
  /* fppowtf32.vhdl:4886:44  */
  assign n4253 = fixrealkcm_freq500_uid89_t1[1]; // extract
  /* fppowtf32.vhdl:4887:44  */
  assign n4254 = fixrealkcm_freq500_uid89_t1[2]; // extract
  /* fppowtf32.vhdl:4888:44  */
  assign n4255 = fixrealkcm_freq500_uid89_t1[3]; // extract
  /* fppowtf32.vhdl:4889:44  */
  assign n4256 = fixrealkcm_freq500_uid89_t1[4]; // extract
  /* fppowtf32.vhdl:4890:44  */
  assign n4257 = fixrealkcm_freq500_uid89_t1[5]; // extract
  /* fppowtf32.vhdl:4891:44  */
  assign n4258 = fixrealkcm_freq500_uid89_t1[6]; // extract
  /* fppowtf32.vhdl:4892:44  */
  assign n4259 = fixrealkcm_freq500_uid89_t1[7]; // extract
  /* fppowtf32.vhdl:4893:44  */
  assign n4260 = fixrealkcm_freq500_uid89_t1[8]; // extract
  /* fppowtf32.vhdl:4894:44  */
  assign n4261 = fixrealkcm_freq500_uid89_t1[9]; // extract
  /* fppowtf32.vhdl:4895:45  */
  assign n4262 = fixrealkcm_freq500_uid89_t1[10]; // extract
  /* fppowtf32.vhdl:4896:45  */
  assign n4263 = fixrealkcm_freq500_uid89_t1[11]; // extract
  /* fppowtf32.vhdl:4897:45  */
  assign n4264 = fixrealkcm_freq500_uid89_t1[12]; // extract
  /* fppowtf32.vhdl:4898:45  */
  assign n4265 = fixrealkcm_freq500_uid89_t1[13]; // extract
  /* fppowtf32.vhdl:4899:45  */
  assign n4266 = fixrealkcm_freq500_uid89_t1[14]; // extract
  /* fppowtf32.vhdl:4900:45  */
  assign n4267 = fixrealkcm_freq500_uid89_t1[15]; // extract
  /* fppowtf32.vhdl:4906:48  */
  assign n4269 = {bh90_w20_0, bh90_w19_0};
  /* fppowtf32.vhdl:4906:61  */
  assign n4270 = {n4269, bh90_w18_0};
  /* fppowtf32.vhdl:4906:74  */
  assign n4271 = {n4270, bh90_w17_0};
  /* fppowtf32.vhdl:4906:87  */
  assign n4272 = {n4271, bh90_w16_0};
  /* fppowtf32.vhdl:4906:100  */
  assign n4273 = {n4272, bh90_w15_0};
  /* fppowtf32.vhdl:4906:113  */
  assign n4274 = {n4273, bh90_w14_0};
  /* fppowtf32.vhdl:4906:126  */
  assign n4275 = {n4274, bh90_w13_0};
  /* fppowtf32.vhdl:4906:139  */
  assign n4276 = {n4275, bh90_w12_0};
  /* fppowtf32.vhdl:4906:152  */
  assign n4277 = {n4276, bh90_w11_0};
  /* fppowtf32.vhdl:4906:165  */
  assign n4278 = {n4277, bh90_w10_0};
  /* fppowtf32.vhdl:4906:178  */
  assign n4279 = {n4278, bh90_w9_0};
  /* fppowtf32.vhdl:4906:190  */
  assign n4280 = {n4279, bh90_w8_0};
  /* fppowtf32.vhdl:4906:202  */
  assign n4281 = {n4280, bh90_w7_0};
  /* fppowtf32.vhdl:4906:214  */
  assign n4282 = {n4281, bh90_w6_0};
  /* fppowtf32.vhdl:4906:226  */
  assign n4283 = {n4282, bh90_w5_0};
  /* fppowtf32.vhdl:4906:238  */
  assign n4284 = {n4283, bh90_w4_0};
  /* fppowtf32.vhdl:4906:250  */
  assign n4285 = {n4284, bh90_w3_0};
  /* fppowtf32.vhdl:4906:262  */
  assign n4286 = {n4285, bh90_w2_0};
  /* fppowtf32.vhdl:4906:274  */
  assign n4287 = {n4286, bh90_w1_0};
  /* fppowtf32.vhdl:4906:286  */
  assign n4288 = {n4287, bh90_w0_0};
  /* fppowtf32.vhdl:4907:60  */
  assign n4290 = {5'b00000, bh90_w15_1};
  /* fppowtf32.vhdl:4907:73  */
  assign n4291 = {n4290, bh90_w14_1};
  /* fppowtf32.vhdl:4907:86  */
  assign n4292 = {n4291, bh90_w13_1};
  /* fppowtf32.vhdl:4907:99  */
  assign n4293 = {n4292, bh90_w12_1};
  /* fppowtf32.vhdl:4907:112  */
  assign n4294 = {n4293, bh90_w11_1};
  /* fppowtf32.vhdl:4907:125  */
  assign n4295 = {n4294, bh90_w10_1};
  /* fppowtf32.vhdl:4907:138  */
  assign n4296 = {n4295, bh90_w9_1};
  /* fppowtf32.vhdl:4907:150  */
  assign n4297 = {n4296, bh90_w8_1};
  /* fppowtf32.vhdl:4907:162  */
  assign n4298 = {n4297, bh90_w7_1};
  /* fppowtf32.vhdl:4907:174  */
  assign n4299 = {n4298, bh90_w6_1};
  /* fppowtf32.vhdl:4907:186  */
  assign n4300 = {n4299, bh90_w5_1};
  /* fppowtf32.vhdl:4907:198  */
  assign n4301 = {n4300, bh90_w4_1};
  /* fppowtf32.vhdl:4907:210  */
  assign n4302 = {n4301, bh90_w3_1};
  /* fppowtf32.vhdl:4907:222  */
  assign n4303 = {n4302, bh90_w2_1};
  /* fppowtf32.vhdl:4907:234  */
  assign n4304 = {n4303, bh90_w1_1};
  /* fppowtf32.vhdl:4907:246  */
  assign n4305 = {n4304, bh90_w0_1};
  /* fppowtf32.vhdl:4910:4  */
  intadder_21_freq500_uid99 bitheapfinaladd_bh90 (
    .clk(clk),
    .x(bitheapfinaladd_bh90_in0),
    .y(bitheapfinaladd_bh90_in1),
    .cin(bitheapfinaladd_bh90_cin),
    .r(bitheapfinaladd_bh90_n4307));
endmodule

module fixrealkcm_freq500_uid77
  (input  clk,
   input  [9:0] x,
   output [7:0] r);
  wire [4:0] fixrealkcm_freq500_uid77_a0;
  wire [11:0] fixrealkcm_freq500_uid77_t0;
  wire [11:0] fixrealkcm_freq500_uid77_t0_copy81;
  wire bh78_w0_0;
  wire bh78_w1_0;
  wire bh78_w2_0;
  wire bh78_w3_0;
  wire bh78_w4_0;
  wire bh78_w5_0;
  wire bh78_w6_0;
  wire bh78_w7_0;
  wire bh78_w8_0;
  wire bh78_w9_0;
  wire bh78_w10_0;
  wire bh78_w11_0;
  wire [4:0] fixrealkcm_freq500_uid77_a1;
  wire [6:0] fixrealkcm_freq500_uid77_t1;
  wire [6:0] fixrealkcm_freq500_uid77_t1_copy84;
  wire bh78_w0_1;
  wire bh78_w1_1;
  wire bh78_w2_1;
  wire bh78_w3_1;
  wire bh78_w4_1;
  wire bh78_w5_1;
  wire bh78_w6_1;
  wire [11:0] bitheapfinaladd_bh78_in0;
  wire [11:0] bitheapfinaladd_bh78_in1;
  wire bitheapfinaladd_bh78_cin;
  wire [11:0] bitheapfinaladd_bh78_out;
  wire [11:0] bitheapresult_bh78;
  wire [11:0] outres;
  wire [4:0] n4170;
  wire [11:0] fixrealkcm_freq500_uid77_table0_n4171;
  wire n4174;
  wire n4175;
  wire n4176;
  wire n4177;
  wire n4178;
  wire n4179;
  wire n4180;
  wire n4181;
  wire n4182;
  wire n4183;
  wire n4184;
  wire n4185;
  wire [4:0] n4186;
  wire [6:0] fixrealkcm_freq500_uid77_table1_n4187;
  wire n4190;
  wire n4191;
  wire n4192;
  wire n4193;
  wire n4194;
  wire n4195;
  wire n4196;
  wire [1:0] n4198;
  wire [2:0] n4199;
  wire [3:0] n4200;
  wire [4:0] n4201;
  wire [5:0] n4202;
  wire [6:0] n4203;
  wire [7:0] n4204;
  wire [8:0] n4205;
  wire [9:0] n4206;
  wire [10:0] n4207;
  wire [11:0] n4208;
  wire [5:0] n4210;
  wire [6:0] n4211;
  wire [7:0] n4212;
  wire [8:0] n4213;
  wire [9:0] n4214;
  wire [10:0] n4215;
  wire [11:0] n4216;
  wire [11:0] bitheapfinaladd_bh78_n4218;
  wire [7:0] n4221;
  assign r = n4221; //(module output)
  /* fppowtf32.vhdl:4524:8  */
  assign fixrealkcm_freq500_uid77_a0 = n4170; // (signal)
  /* fppowtf32.vhdl:4526:8  */
  assign fixrealkcm_freq500_uid77_t0 = fixrealkcm_freq500_uid77_t0_copy81; // (signal)
  /* fppowtf32.vhdl:4528:8  */
  assign fixrealkcm_freq500_uid77_t0_copy81 = fixrealkcm_freq500_uid77_table0_n4171; // (signal)
  /* fppowtf32.vhdl:4530:8  */
  assign bh78_w0_0 = n4174; // (signal)
  /* fppowtf32.vhdl:4532:8  */
  assign bh78_w1_0 = n4175; // (signal)
  /* fppowtf32.vhdl:4534:8  */
  assign bh78_w2_0 = n4176; // (signal)
  /* fppowtf32.vhdl:4536:8  */
  assign bh78_w3_0 = n4177; // (signal)
  /* fppowtf32.vhdl:4538:8  */
  assign bh78_w4_0 = n4178; // (signal)
  /* fppowtf32.vhdl:4540:8  */
  assign bh78_w5_0 = n4179; // (signal)
  /* fppowtf32.vhdl:4542:8  */
  assign bh78_w6_0 = n4180; // (signal)
  /* fppowtf32.vhdl:4544:8  */
  assign bh78_w7_0 = n4181; // (signal)
  /* fppowtf32.vhdl:4546:8  */
  assign bh78_w8_0 = n4182; // (signal)
  /* fppowtf32.vhdl:4548:8  */
  assign bh78_w9_0 = n4183; // (signal)
  /* fppowtf32.vhdl:4550:8  */
  assign bh78_w10_0 = n4184; // (signal)
  /* fppowtf32.vhdl:4622:35  */
  assign bh78_w11_0 = n4185; // (signal)
  /* fppowtf32.vhdl:4554:8  */
  assign fixrealkcm_freq500_uid77_a1 = n4186; // (signal)
  /* fppowtf32.vhdl:4556:8  */
  assign fixrealkcm_freq500_uid77_t1 = fixrealkcm_freq500_uid77_t1_copy84; // (signal)
  /* fppowtf32.vhdl:4558:8  */
  assign fixrealkcm_freq500_uid77_t1_copy84 = fixrealkcm_freq500_uid77_table1_n4187; // (signal)
  /* fppowtf32.vhdl:4560:8  */
  assign bh78_w0_1 = n4190; // (signal)
  /* fppowtf32.vhdl:4562:8  */
  assign bh78_w1_1 = n4191; // (signal)
  /* fppowtf32.vhdl:4564:8  */
  assign bh78_w2_1 = n4192; // (signal)
  /* fppowtf32.vhdl:4566:8  */
  assign bh78_w3_1 = n4193; // (signal)
  /* fppowtf32.vhdl:4568:8  */
  assign bh78_w4_1 = n4194; // (signal)
  /* fppowtf32.vhdl:4570:8  */
  assign bh78_w5_1 = n4195; // (signal)
  /* fppowtf32.vhdl:4572:8  */
  assign bh78_w6_1 = n4196; // (signal)
  /* fppowtf32.vhdl:4574:8  */
  assign bitheapfinaladd_bh78_in0 = n4208; // (signal)
  /* fppowtf32.vhdl:4576:8  */
  assign bitheapfinaladd_bh78_in1 = n4216; // (signal)
  /* fppowtf32.vhdl:4578:8  */
  assign bitheapfinaladd_bh78_cin = 1'b0; // (signal)
  /* fppowtf32.vhdl:4580:8  */
  assign bitheapfinaladd_bh78_out = bitheapfinaladd_bh78_n4218; // (signal)
  /* fppowtf32.vhdl:4582:8  */
  assign bitheapresult_bh78 = bitheapfinaladd_bh78_out; // (signal)
  /* fppowtf32.vhdl:4584:8  */
  assign outres = bitheapresult_bh78; // (signal)
  /* fppowtf32.vhdl:4588:36  */
  assign n4170 = x[9:5]; // extract
  /* fppowtf32.vhdl:4589:4  */
  fixrealkcm_freq500_uid77_t0_freq500_uid80 fixrealkcm_freq500_uid77_table0 (
    .x(fixrealkcm_freq500_uid77_a0),
    .y(fixrealkcm_freq500_uid77_table0_n4171));
  /* fppowtf32.vhdl:4593:44  */
  assign n4174 = fixrealkcm_freq500_uid77_t0[0]; // extract
  /* fppowtf32.vhdl:4594:44  */
  assign n4175 = fixrealkcm_freq500_uid77_t0[1]; // extract
  /* fppowtf32.vhdl:4595:44  */
  assign n4176 = fixrealkcm_freq500_uid77_t0[2]; // extract
  /* fppowtf32.vhdl:4596:44  */
  assign n4177 = fixrealkcm_freq500_uid77_t0[3]; // extract
  /* fppowtf32.vhdl:4597:44  */
  assign n4178 = fixrealkcm_freq500_uid77_t0[4]; // extract
  /* fppowtf32.vhdl:4598:44  */
  assign n4179 = fixrealkcm_freq500_uid77_t0[5]; // extract
  /* fppowtf32.vhdl:4599:44  */
  assign n4180 = fixrealkcm_freq500_uid77_t0[6]; // extract
  /* fppowtf32.vhdl:4600:44  */
  assign n4181 = fixrealkcm_freq500_uid77_t0[7]; // extract
  /* fppowtf32.vhdl:4601:44  */
  assign n4182 = fixrealkcm_freq500_uid77_t0[8]; // extract
  /* fppowtf32.vhdl:4602:44  */
  assign n4183 = fixrealkcm_freq500_uid77_t0[9]; // extract
  /* fppowtf32.vhdl:4603:45  */
  assign n4184 = fixrealkcm_freq500_uid77_t0[10]; // extract
  /* fppowtf32.vhdl:4604:45  */
  assign n4185 = fixrealkcm_freq500_uid77_t0[11]; // extract
  /* fppowtf32.vhdl:4605:36  */
  assign n4186 = x[4:0]; // extract
  /* fppowtf32.vhdl:4606:4  */
  fixrealkcm_freq500_uid77_t1_freq500_uid83 fixrealkcm_freq500_uid77_table1 (
    .x(fixrealkcm_freq500_uid77_a1),
    .y(fixrealkcm_freq500_uid77_table1_n4187));
  /* fppowtf32.vhdl:4610:44  */
  assign n4190 = fixrealkcm_freq500_uid77_t1[0]; // extract
  /* fppowtf32.vhdl:4611:44  */
  assign n4191 = fixrealkcm_freq500_uid77_t1[1]; // extract
  /* fppowtf32.vhdl:4612:44  */
  assign n4192 = fixrealkcm_freq500_uid77_t1[2]; // extract
  /* fppowtf32.vhdl:4613:44  */
  assign n4193 = fixrealkcm_freq500_uid77_t1[3]; // extract
  /* fppowtf32.vhdl:4614:44  */
  assign n4194 = fixrealkcm_freq500_uid77_t1[4]; // extract
  /* fppowtf32.vhdl:4615:44  */
  assign n4195 = fixrealkcm_freq500_uid77_t1[5]; // extract
  /* fppowtf32.vhdl:4616:44  */
  assign n4196 = fixrealkcm_freq500_uid77_t1[6]; // extract
  /* fppowtf32.vhdl:4622:48  */
  assign n4198 = {bh78_w11_0, bh78_w10_0};
  /* fppowtf32.vhdl:4622:61  */
  assign n4199 = {n4198, bh78_w9_0};
  /* fppowtf32.vhdl:4622:73  */
  assign n4200 = {n4199, bh78_w8_0};
  /* fppowtf32.vhdl:4622:85  */
  assign n4201 = {n4200, bh78_w7_0};
  /* fppowtf32.vhdl:4622:97  */
  assign n4202 = {n4201, bh78_w6_0};
  /* fppowtf32.vhdl:4622:109  */
  assign n4203 = {n4202, bh78_w5_0};
  /* fppowtf32.vhdl:4622:121  */
  assign n4204 = {n4203, bh78_w4_0};
  /* fppowtf32.vhdl:4622:133  */
  assign n4205 = {n4204, bh78_w3_0};
  /* fppowtf32.vhdl:4622:145  */
  assign n4206 = {n4205, bh78_w2_0};
  /* fppowtf32.vhdl:4622:157  */
  assign n4207 = {n4206, bh78_w1_0};
  /* fppowtf32.vhdl:4622:169  */
  assign n4208 = {n4207, bh78_w0_0};
  /* fppowtf32.vhdl:4623:60  */
  assign n4210 = {5'b00000, bh78_w6_1};
  /* fppowtf32.vhdl:4623:72  */
  assign n4211 = {n4210, bh78_w5_1};
  /* fppowtf32.vhdl:4623:84  */
  assign n4212 = {n4211, bh78_w4_1};
  /* fppowtf32.vhdl:4623:96  */
  assign n4213 = {n4212, bh78_w3_1};
  /* fppowtf32.vhdl:4623:108  */
  assign n4214 = {n4213, bh78_w2_1};
  /* fppowtf32.vhdl:4623:120  */
  assign n4215 = {n4214, bh78_w1_1};
  /* fppowtf32.vhdl:4623:132  */
  assign n4216 = {n4215, bh78_w0_1};
  /* fppowtf32.vhdl:4626:4  */
  intadder_12_freq500_uid87 bitheapfinaladd_bh78 (
    .clk(clk),
    .x(bitheapfinaladd_bh78_in0),
    .y(bitheapfinaladd_bh78_in1),
    .cin(bitheapfinaladd_bh78_cin),
    .r(bitheapfinaladd_bh78_n4218));
  /* fppowtf32.vhdl:4634:15  */
  assign n4221 = outres[11:4]; // extract
endmodule

module intadder_32_freq500_uid49
  (input  clk,
   input  [31:0] x,
   input  [31:0] y,
   input  cin,
   output [31:0] r);
  wire [31:0] rtmp;
  wire cin_d1;
  wire [31:0] n4165;
  wire [31:0] n4166;
  wire [31:0] n4167;
  reg n4168;
  assign r = rtmp; //(module output)
  /* fppowtf32.vhdl:2797:8  */
  assign rtmp = n4167; // (signal)
  /* fppowtf32.vhdl:2799:8  */
  assign cin_d1 = n4168; // (signal)
  /* fppowtf32.vhdl:2808:14  */
  assign n4165 = x + y;
  /* fppowtf32.vhdl:2808:18  */
  assign n4166 = {31'b0, cin_d1};  //  uext
  /* fppowtf32.vhdl:2808:18  */
  assign n4167 = n4165 + n4166;
  /* fppowtf32.vhdl:2804:10  */
  always @(posedge clk)
    n4168 <= cin;
endmodule

module fixrealkcm_freq500_uid39_t1_freq500_uid45
  (input  [2:0] x,
   output [26:0] y);
  wire [26:0] y0;
  wire [26:0] y1;
  wire n4134;
  wire n4137;
  wire n4140;
  wire n4143;
  wire n4146;
  wire n4149;
  wire n4152;
  wire n4155;
  wire [7:0] n4157;
  reg [26:0] n4158;
  assign y = y1; //(module output)
  /* fppowtf32.vhdl:798:8  */
  assign y0 = n4158; // (signal)
  /* fppowtf32.vhdl:800:8  */
  assign y1 = y0; // (signal)
  /* fppowtf32.vhdl:804:37  */
  assign n4134 = x == 3'b000;
  /* fppowtf32.vhdl:805:37  */
  assign n4137 = x == 3'b001;
  /* fppowtf32.vhdl:806:37  */
  assign n4140 = x == 3'b010;
  /* fppowtf32.vhdl:807:37  */
  assign n4143 = x == 3'b011;
  /* fppowtf32.vhdl:808:37  */
  assign n4146 = x == 3'b100;
  /* fppowtf32.vhdl:809:37  */
  assign n4149 = x == 3'b101;
  /* fppowtf32.vhdl:810:37  */
  assign n4152 = x == 3'b110;
  /* fppowtf32.vhdl:811:37  */
  assign n4155 = x == 3'b111;
  assign n4157 = {n4155, n4152, n4149, n4146, n4143, n4140, n4137, n4134};
  /* fppowtf32.vhdl:803:4  */
  always @*
    case (n4157)
      8'b10000000: n4158 = 27'b100110110100001111010101000;
      8'b01000000: n4158 = 27'b100001010001010110010010000;
      8'b00100000: n4158 = 27'b011011101110011101001111000;
      8'b00010000: n4158 = 27'b010110001011100100001100000;
      8'b00001000: n4158 = 27'b010000101000101011001001000;
      8'b00000100: n4158 = 27'b001011000101110010000110000;
      8'b00000010: n4158 = 27'b000101100010111001000011000;
      8'b00000001: n4158 = 27'b000000000000000000000000000;
      default: n4158 = 27'bX;
    endcase
endmodule

module fixrealkcm_freq500_uid39_t0_freq500_uid42
  (input  [4:0] x,
   output [31:0] y);
  wire [31:0] y0;
  wire [31:0] y1;
  wire n4034;
  wire n4037;
  wire n4040;
  wire n4043;
  wire n4046;
  wire n4049;
  wire n4052;
  wire n4055;
  wire n4058;
  wire n4061;
  wire n4064;
  wire n4067;
  wire n4070;
  wire n4073;
  wire n4076;
  wire n4079;
  wire n4082;
  wire n4085;
  wire n4088;
  wire n4091;
  wire n4094;
  wire n4097;
  wire n4100;
  wire n4103;
  wire n4106;
  wire n4109;
  wire n4112;
  wire n4115;
  wire n4118;
  wire n4121;
  wire n4124;
  wire n4127;
  wire [31:0] n4129;
  reg [31:0] n4130;
  assign y = y1; //(module output)
  /* fppowtf32.vhdl:726:8  */
  assign y0 = n4130; // (signal)
  /* fppowtf32.vhdl:728:8  */
  assign y1 = y0; // (signal)
  /* fppowtf32.vhdl:732:42  */
  assign n4034 = x == 5'b00000;
  /* fppowtf32.vhdl:733:42  */
  assign n4037 = x == 5'b00001;
  /* fppowtf32.vhdl:734:42  */
  assign n4040 = x == 5'b00010;
  /* fppowtf32.vhdl:735:42  */
  assign n4043 = x == 5'b00011;
  /* fppowtf32.vhdl:736:42  */
  assign n4046 = x == 5'b00100;
  /* fppowtf32.vhdl:737:42  */
  assign n4049 = x == 5'b00101;
  /* fppowtf32.vhdl:738:42  */
  assign n4052 = x == 5'b00110;
  /* fppowtf32.vhdl:739:42  */
  assign n4055 = x == 5'b00111;
  /* fppowtf32.vhdl:740:42  */
  assign n4058 = x == 5'b01000;
  /* fppowtf32.vhdl:741:42  */
  assign n4061 = x == 5'b01001;
  /* fppowtf32.vhdl:742:42  */
  assign n4064 = x == 5'b01010;
  /* fppowtf32.vhdl:743:42  */
  assign n4067 = x == 5'b01011;
  /* fppowtf32.vhdl:744:42  */
  assign n4070 = x == 5'b01100;
  /* fppowtf32.vhdl:745:42  */
  assign n4073 = x == 5'b01101;
  /* fppowtf32.vhdl:746:42  */
  assign n4076 = x == 5'b01110;
  /* fppowtf32.vhdl:747:42  */
  assign n4079 = x == 5'b01111;
  /* fppowtf32.vhdl:748:42  */
  assign n4082 = x == 5'b10000;
  /* fppowtf32.vhdl:749:42  */
  assign n4085 = x == 5'b10001;
  /* fppowtf32.vhdl:750:42  */
  assign n4088 = x == 5'b10010;
  /* fppowtf32.vhdl:751:42  */
  assign n4091 = x == 5'b10011;
  /* fppowtf32.vhdl:752:42  */
  assign n4094 = x == 5'b10100;
  /* fppowtf32.vhdl:753:42  */
  assign n4097 = x == 5'b10101;
  /* fppowtf32.vhdl:754:42  */
  assign n4100 = x == 5'b10110;
  /* fppowtf32.vhdl:755:42  */
  assign n4103 = x == 5'b10111;
  /* fppowtf32.vhdl:756:42  */
  assign n4106 = x == 5'b11000;
  /* fppowtf32.vhdl:757:42  */
  assign n4109 = x == 5'b11001;
  /* fppowtf32.vhdl:758:42  */
  assign n4112 = x == 5'b11010;
  /* fppowtf32.vhdl:759:42  */
  assign n4115 = x == 5'b11011;
  /* fppowtf32.vhdl:760:42  */
  assign n4118 = x == 5'b11100;
  /* fppowtf32.vhdl:761:42  */
  assign n4121 = x == 5'b11101;
  /* fppowtf32.vhdl:762:42  */
  assign n4124 = x == 5'b11110;
  /* fppowtf32.vhdl:763:42  */
  assign n4127 = x == 5'b11111;
  assign n4129 = {n4127, n4124, n4121, n4118, n4115, n4112, n4109, n4106, n4103, n4100, n4097, n4094, n4091, n4088, n4085, n4082, n4079, n4076, n4073, n4070, n4067, n4064, n4061, n4058, n4055, n4052, n4049, n4046, n4043, n4040, n4037, n4034};
  /* fppowtf32.vhdl:731:4  */
  always @*
    case (n4129)
      32'b10000000000000000000000000000000: n4130 = 32'b10101011111001101000011100111000;
      32'b01000000000000000000000000000000: n4130 = 32'b10100110010110101111011001111000;
      32'b00100000000000000000000000000000: n4130 = 32'b10100000110011110110010110111001;
      32'b00010000000000000000000000000000: n4130 = 32'b10011011010000111101010011111001;
      32'b00001000000000000000000000000000: n4130 = 32'b10010101101110000100010000111001;
      32'b00000100000000000000000000000000: n4130 = 32'b10010000001011001011001101111001;
      32'b00000010000000000000000000000000: n4130 = 32'b10001010101000010010001010111010;
      32'b00000001000000000000000000000000: n4130 = 32'b10000101000101011001000111111010;
      32'b00000000100000000000000000000000: n4130 = 32'b01111111100010100000000100111010;
      32'b00000000010000000000000000000000: n4130 = 32'b01111001111111100111000001111010;
      32'b00000000001000000000000000000000: n4130 = 32'b01110100011100101101111110111011;
      32'b00000000000100000000000000000000: n4130 = 32'b01101110111001110100111011111011;
      32'b00000000000010000000000000000000: n4130 = 32'b01101001010110111011111000111011;
      32'b00000000000001000000000000000000: n4130 = 32'b01100011110100000010110101111011;
      32'b00000000000000100000000000000000: n4130 = 32'b01011110010001001001110010111100;
      32'b00000000000000010000000000000000: n4130 = 32'b01011000101110010000101111111100;
      32'b00000000000000001000000000000000: n4130 = 32'b01010011001011010111101100111100;
      32'b00000000000000000100000000000000: n4130 = 32'b01001101101000011110101001111100;
      32'b00000000000000000010000000000000: n4130 = 32'b01001000000101100101100110111101;
      32'b00000000000000000001000000000000: n4130 = 32'b01000010100010101100100011111101;
      32'b00000000000000000000100000000000: n4130 = 32'b00111100111111110011100000111101;
      32'b00000000000000000000010000000000: n4130 = 32'b00110111011100111010011101111101;
      32'b00000000000000000000001000000000: n4130 = 32'b00110001111010000001011010111110;
      32'b00000000000000000000000100000000: n4130 = 32'b00101100010111001000010111111110;
      32'b00000000000000000000000010000000: n4130 = 32'b00100110110100001111010100111110;
      32'b00000000000000000000000001000000: n4130 = 32'b00100001010001010110010001111110;
      32'b00000000000000000000000000100000: n4130 = 32'b00011011101110011101001110111111;
      32'b00000000000000000000000000010000: n4130 = 32'b00010110001011100100001011111111;
      32'b00000000000000000000000000001000: n4130 = 32'b00010000101000101011001000111111;
      32'b00000000000000000000000000000100: n4130 = 32'b00001011000101110010000101111111;
      32'b00000000000000000000000000000010: n4130 = 32'b00000101100010111001000011000000;
      32'b00000000000000000000000000000001: n4130 = 32'b00000000000000000000000000000000;
      default: n4130 = 32'bX;
    endcase
endmodule

module intadder_20_freq500_uid121
  (input  clk,
   input  [19:0] x,
   input  [19:0] y,
   input  cin,
   output [19:0] r);
  wire [19:0] rtmp;
  wire [19:0] x_d1;
  wire [19:0] y_d1;
  wire cin_d1;
  wire cin_d2;
  wire cin_d3;
  wire cin_d4;
  wire cin_d5;
  wire cin_d6;
  wire cin_d7;
  wire cin_d8;
  wire cin_d9;
  wire cin_d10;
  wire cin_d11;
  wire cin_d12;
  wire cin_d13;
  wire cin_d14;
  wire cin_d15;
  wire cin_d16;
  wire cin_d17;
  wire cin_d18;
  wire cin_d19;
  wire cin_d20;
  wire [19:0] n4006;
  wire [19:0] n4007;
  wire [19:0] n4008;
  reg [19:0] n4009;
  reg [19:0] n4010;
  reg n4011;
  reg n4012;
  reg n4013;
  reg n4014;
  reg n4015;
  reg n4016;
  reg n4017;
  reg n4018;
  reg n4019;
  reg n4020;
  reg n4021;
  reg n4022;
  reg n4023;
  reg n4024;
  reg n4025;
  reg n4026;
  reg n4027;
  reg n4028;
  reg n4029;
  reg n4030;
  assign r = rtmp; //(module output)
  /* fppowtf32.vhdl:5436:8  */
  assign rtmp = n4008; // (signal)
  /* fppowtf32.vhdl:5438:8  */
  assign x_d1 = n4009; // (signal)
  /* fppowtf32.vhdl:5440:8  */
  assign y_d1 = n4010; // (signal)
  /* fppowtf32.vhdl:5442:8  */
  assign cin_d1 = n4011; // (signal)
  /* fppowtf32.vhdl:5442:16  */
  assign cin_d2 = n4012; // (signal)
  /* fppowtf32.vhdl:5442:24  */
  assign cin_d3 = n4013; // (signal)
  /* fppowtf32.vhdl:5442:32  */
  assign cin_d4 = n4014; // (signal)
  /* fppowtf32.vhdl:5442:40  */
  assign cin_d5 = n4015; // (signal)
  /* fppowtf32.vhdl:5442:48  */
  assign cin_d6 = n4016; // (signal)
  /* fppowtf32.vhdl:5442:56  */
  assign cin_d7 = n4017; // (signal)
  /* fppowtf32.vhdl:5442:64  */
  assign cin_d8 = n4018; // (signal)
  /* fppowtf32.vhdl:5442:72  */
  assign cin_d9 = n4019; // (signal)
  /* fppowtf32.vhdl:5442:80  */
  assign cin_d10 = n4020; // (signal)
  /* fppowtf32.vhdl:5442:89  */
  assign cin_d11 = n4021; // (signal)
  /* fppowtf32.vhdl:5442:98  */
  assign cin_d12 = n4022; // (signal)
  /* fppowtf32.vhdl:5442:107  */
  assign cin_d13 = n4023; // (signal)
  /* fppowtf32.vhdl:5442:116  */
  assign cin_d14 = n4024; // (signal)
  /* fppowtf32.vhdl:5442:125  */
  assign cin_d15 = n4025; // (signal)
  /* fppowtf32.vhdl:5442:134  */
  assign cin_d16 = n4026; // (signal)
  /* fppowtf32.vhdl:5442:143  */
  assign cin_d17 = n4027; // (signal)
  /* fppowtf32.vhdl:5442:152  */
  assign cin_d18 = n4028; // (signal)
  /* fppowtf32.vhdl:5442:161  */
  assign cin_d19 = n4029; // (signal)
  /* fppowtf32.vhdl:5442:170  */
  assign cin_d20 = n4030; // (signal)
  /* fppowtf32.vhdl:5472:17  */
  assign n4006 = x_d1 + y_d1;
  /* fppowtf32.vhdl:5472:24  */
  assign n4007 = {19'b0, cin_d20};  //  uext
  /* fppowtf32.vhdl:5472:24  */
  assign n4008 = n4006 + n4007;
  /* fppowtf32.vhdl:5447:10  */
  always @(posedge clk)
    n4009 <= x;
  /* fppowtf32.vhdl:5447:10  */
  always @(posedge clk)
    n4010 <= y;
  /* fppowtf32.vhdl:5447:10  */
  always @(posedge clk)
    n4011 <= cin;
  /* fppowtf32.vhdl:5447:10  */
  always @(posedge clk)
    n4012 <= cin_d1;
  /* fppowtf32.vhdl:5447:10  */
  always @(posedge clk)
    n4013 <= cin_d2;
  /* fppowtf32.vhdl:5447:10  */
  always @(posedge clk)
    n4014 <= cin_d3;
  /* fppowtf32.vhdl:5447:10  */
  always @(posedge clk)
    n4015 <= cin_d4;
  /* fppowtf32.vhdl:5447:10  */
  always @(posedge clk)
    n4016 <= cin_d5;
  /* fppowtf32.vhdl:5447:10  */
  always @(posedge clk)
    n4017 <= cin_d6;
  /* fppowtf32.vhdl:5447:10  */
  always @(posedge clk)
    n4018 <= cin_d7;
  /* fppowtf32.vhdl:5447:10  */
  always @(posedge clk)
    n4019 <= cin_d8;
  /* fppowtf32.vhdl:5447:10  */
  always @(posedge clk)
    n4020 <= cin_d9;
  /* fppowtf32.vhdl:5447:10  */
  always @(posedge clk)
    n4021 <= cin_d10;
  /* fppowtf32.vhdl:5447:10  */
  always @(posedge clk)
    n4022 <= cin_d11;
  /* fppowtf32.vhdl:5447:10  */
  always @(posedge clk)
    n4023 <= cin_d12;
  /* fppowtf32.vhdl:5447:10  */
  always @(posedge clk)
    n4024 <= cin_d13;
  /* fppowtf32.vhdl:5447:10  */
  always @(posedge clk)
    n4025 <= cin_d14;
  /* fppowtf32.vhdl:5447:10  */
  always @(posedge clk)
    n4026 <= cin_d15;
  /* fppowtf32.vhdl:5447:10  */
  always @(posedge clk)
    n4027 <= cin_d16;
  /* fppowtf32.vhdl:5447:10  */
  always @(posedge clk)
    n4028 <= cin_d17;
  /* fppowtf32.vhdl:5447:10  */
  always @(posedge clk)
    n4029 <= cin_d18;
  /* fppowtf32.vhdl:5447:10  */
  always @(posedge clk)
    n4030 <= cin_d19;
endmodule

module exp_8_10_freq500_uid75
  (input  clk,
   input  [19:0] ufixx_i,
   input  xsign,
   output [13:0] expy,
   output [8:0] k);
  wire [19:0] ufixx;
  wire [9:0] xmulin;
  wire [7:0] absk;
  wire [7:0] absk_d1;
  wire [8:0] minusabsk;
  wire [20:0] absklog2;
  wire [12:0] subop1;
  wire [12:0] subop2;
  wire [12:0] y;
  wire [9:0] a;
  wire [2:0] z;
  wire [13:0] expa;
  wire [13:0] expa_copy105;
  wire [2:0] expzm1_p;
  wire [2:0] expzm1_p_copy108;
  wire [3:0] expzm1;
  wire [3:0] expa_t;
  wire [3:0] exparounded0;
  wire [2:0] exparounded;
  wire [4:0] lowerproduct;
  wire [13:0] extendedlowerproduct;
  wire xsign_d1;
  wire xsign_d2;
  wire xsign_d3;
  wire xsign_d4;
  wire [9:0] n3921;
  wire [7:0] mulinvlog2_n3922;
  wire [8:0] n3926;
  wire [8:0] n3928;
  wire [8:0] n3929;
  wire [8:0] n3931;
  wire [20:0] mullog2_n3932;
  wire [12:0] n3935;
  wire n3936;
  wire [12:0] n3937;
  wire [12:0] n3938;
  wire [12:0] n3939;
  wire [12:0] n3940;
  wire [12:0] n3941;
  wire [12:0] n3942;
  wire [12:0] n3943;
  localparam n3944 = 1'b1;
  wire [12:0] theyadder_n3945;
  wire [9:0] n3948;
  wire [2:0] n3949;
  wire [13:0] expatable_n3950;
  wire [2:0] expzm1table_n3953;
  wire [3:0] n3957;
  wire [3:0] n3958;
  localparam [3:0] n3959 = 4'b0000;
  localparam n3960 = 1'b1;
  wire [3:0] adder_exparounded0_n3961;
  wire [2:0] n3964;
  wire [4:0] thelowerproduct_n3965;
  wire [13:0] n3969;
  localparam n3970 = 1'b0;
  wire [13:0] thefinaladder_n3971;
  reg [7:0] n3974;
  reg n3975;
  reg n3976;
  reg n3977;
  reg n3978;
  assign expy = thefinaladder_n3971; //(module output)
  assign k = n3929; //(module output)
  /* fppowtf32.vhdl:5292:8  */
  assign xmulin = n3921; // (signal)
  /* fppowtf32.vhdl:5294:8  */
  assign absk = mulinvlog2_n3922; // (signal)
  /* fppowtf32.vhdl:5294:14  */
  assign absk_d1 = n3974; // (signal)
  /* fppowtf32.vhdl:5296:8  */
  assign minusabsk = n3928; // (signal)
  /* fppowtf32.vhdl:5298:8  */
  assign absklog2 = mullog2_n3932; // (signal)
  /* fppowtf32.vhdl:5300:8  */
  assign subop1 = n3937; // (signal)
  /* fppowtf32.vhdl:5302:8  */
  assign subop2 = n3941; // (signal)
  /* fppowtf32.vhdl:5304:8  */
  assign y = theyadder_n3945; // (signal)
  /* fppowtf32.vhdl:5306:8  */
  assign a = n3948; // (signal)
  /* fppowtf32.vhdl:5308:8  */
  assign z = n3949; // (signal)
  /* fppowtf32.vhdl:5310:8  */
  assign expa = expa_copy105; // (signal)
  /* fppowtf32.vhdl:5312:8  */
  assign expa_copy105 = expatable_n3950; // (signal)
  /* fppowtf32.vhdl:5314:8  */
  assign expzm1_p = expzm1_p_copy108; // (signal)
  /* fppowtf32.vhdl:5316:8  */
  assign expzm1_p_copy108 = expzm1table_n3953; // (signal)
  /* fppowtf32.vhdl:5318:8  */
  assign expzm1 = n3957; // (signal)
  /* fppowtf32.vhdl:5320:8  */
  assign expa_t = n3958; // (signal)
  /* fppowtf32.vhdl:5322:8  */
  assign exparounded0 = adder_exparounded0_n3961; // (signal)
  /* fppowtf32.vhdl:5324:8  */
  assign exparounded = n3964; // (signal)
  /* fppowtf32.vhdl:5326:8  */
  assign lowerproduct = thelowerproduct_n3965; // (signal)
  /* fppowtf32.vhdl:5328:8  */
  assign extendedlowerproduct = n3969; // (signal)
  /* fppowtf32.vhdl:5330:8  */
  assign xsign_d1 = n3975; // (signal)
  /* fppowtf32.vhdl:5330:18  */
  assign xsign_d2 = n3976; // (signal)
  /* fppowtf32.vhdl:5330:28  */
  assign xsign_d3 = n3977; // (signal)
  /* fppowtf32.vhdl:5330:38  */
  assign xsign_d4 = n3978; // (signal)
  /* fppowtf32.vhdl:5348:19  */
  assign n3921 = ufixx[19:10]; // extract
  /* fppowtf32.vhdl:5349:4  */
  fixrealkcm_freq500_uid77 mulinvlog2 (
    .clk(clk),
    .x(xmulin),
    .r(mulinvlog2_n3922));
  /* fppowtf32.vhdl:5353:44  */
  assign n3926 = {1'b0, absk_d1};
  /* fppowtf32.vhdl:5353:37  */
  assign n3928 = 9'b000000000 - n3926;
  /* fppowtf32.vhdl:5354:19  */
  assign n3929 = xsign_d4 ? minusabsk : n3931;
  /* fppowtf32.vhdl:5354:50  */
  assign n3931 = {1'b0, absk_d1};
  /* fppowtf32.vhdl:5355:4  */
  fixrealkcm_freq500_uid89 mullog2 (
    .clk(clk),
    .x(absk),
    .r(mullog2_n3932));
  /* fppowtf32.vhdl:5359:36  */
  assign n3935 = ufixx[12:0]; // extract
  /* fppowtf32.vhdl:5359:64  */
  assign n3936 = ~xsign_d2;
  /* fppowtf32.vhdl:5359:51  */
  assign n3937 = n3936 ? n3935 : n3939;
  /* fppowtf32.vhdl:5359:101  */
  assign n3938 = ufixx[12:0]; // extract
  /* fppowtf32.vhdl:5359:74  */
  assign n3939 = ~n3938;
  /* fppowtf32.vhdl:5360:22  */
  assign n3940 = absklog2[12:0]; // extract
  /* fppowtf32.vhdl:5360:36  */
  assign n3941 = xsign_d4 ? n3940 : n3943;
  /* fppowtf32.vhdl:5360:72  */
  assign n3942 = absklog2[12:0]; // extract
  /* fppowtf32.vhdl:5360:59  */
  assign n3943 = ~n3942;
  /* fppowtf32.vhdl:5361:4  */
  intadder_13_freq500_uid102 theyadder (
    .clk(clk),
    .x(subop1),
    .y(subop2),
    .cin(n3944),
    .r(theyadder_n3945));
  /* fppowtf32.vhdl:5368:10  */
  assign n3948 = y[12:3]; // extract
  /* fppowtf32.vhdl:5369:10  */
  assign n3949 = y[2:0]; // extract
  /* fppowtf32.vhdl:5370:4  */
  fixfunctionbytable_freq500_uid104 expatable (
    .x(a),
    .y(expatable_n3950));
  /* fppowtf32.vhdl:5374:4  */
  fixfunctionbytable_freq500_uid107 expzm1table (
    .x(z),
    .y(expzm1table_n3953));
  /* fppowtf32.vhdl:5378:15  */
  assign n3957 = {1'b0, expzm1_p};
  /* fppowtf32.vhdl:5381:18  */
  assign n3958 = expa[13:10]; // extract
  /* fppowtf32.vhdl:5382:4  */
  intadder_4_freq500_uid112 adder_exparounded0 (
    .clk(clk),
    .x(expa_t),
    .y(n3959),
    .cin(n3960),
    .r(adder_exparounded0_n3961));
  /* fppowtf32.vhdl:5388:31  */
  assign n3964 = exparounded0[3:1]; // extract
  /* fppowtf32.vhdl:5389:4  */
  intmultiplier_3x4_5_freq500_uid114 thelowerproduct (
    .clk(clk),
    .x(exparounded),
    .y(expzm1),
    .r(thelowerproduct_n3965));
  /* fppowtf32.vhdl:5394:50  */
  assign n3969 = {9'b000000000, lowerproduct};
  /* fppowtf32.vhdl:5396:4  */
  intadder_14_freq500_uid118 thefinaladder (
    .clk(clk),
    .x(expa),
    .y(extendedlowerproduct),
    .cin(n3970),
    .r(thefinaladder_n3971));
  /* fppowtf32.vhdl:5339:10  */
  always @(posedge clk)
    n3974 <= absk;
  /* fppowtf32.vhdl:5339:10  */
  always @(posedge clk)
    n3975 <= xsign;
  /* fppowtf32.vhdl:5339:10  */
  always @(posedge clk)
    n3976 <= xsign_d1;
  /* fppowtf32.vhdl:5339:10  */
  always @(posedge clk)
    n3977 <= xsign_d2;
  /* fppowtf32.vhdl:5339:10  */
  always @(posedge clk)
    n3978 <= xsign_d3;
endmodule

module leftshifter22_by_max_19_freq500_uid73
  (input  clk,
   input  [21:0] x,
   input  [4:0] s,
   output [40:0] r);
  wire [4:0] ps;
  wire [4:0] ps_d1;
  wire [21:0] level0;
  wire [21:0] level0_d1;
  wire [22:0] level1;
  wire [22:0] level1_d1;
  wire [24:0] level2;
  wire [28:0] level3;
  wire [36:0] level4;
  wire [52:0] level5;
  wire [22:0] n3877;
  wire n3878;
  wire [22:0] n3879;
  wire [22:0] n3881;
  wire [24:0] n3883;
  wire n3884;
  wire [24:0] n3885;
  wire [24:0] n3887;
  wire [28:0] n3889;
  wire n3890;
  wire [28:0] n3891;
  wire [28:0] n3893;
  wire [36:0] n3895;
  wire n3896;
  wire [36:0] n3897;
  wire [36:0] n3899;
  wire [52:0] n3901;
  wire n3902;
  wire [52:0] n3903;
  wire [52:0] n3905;
  wire [40:0] n3906;
  reg [4:0] n3907;
  reg [21:0] n3908;
  reg [22:0] n3909;
  assign r = n3906; //(module output)
  /* fppowtf32.vhdl:4375:12  */
  assign ps_d1 = n3907; // (signal)
  /* fppowtf32.vhdl:4377:16  */
  assign level0_d1 = n3908; // (signal)
  /* fppowtf32.vhdl:4379:8  */
  assign level1 = n3879; // (signal)
  /* fppowtf32.vhdl:4379:16  */
  assign level1_d1 = n3909; // (signal)
  /* fppowtf32.vhdl:4381:8  */
  assign level2 = n3885; // (signal)
  /* fppowtf32.vhdl:4383:8  */
  assign level3 = n3891; // (signal)
  /* fppowtf32.vhdl:4385:8  */
  assign level4 = n3897; // (signal)
  /* fppowtf32.vhdl:4387:8  */
  assign level5 = n3903; // (signal)
  /* fppowtf32.vhdl:4400:23  */
  assign n3877 = {level0_d1, 1'b0};
  /* fppowtf32.vhdl:4400:52  */
  assign n3878 = ps[0]; // extract
  /* fppowtf32.vhdl:4400:45  */
  assign n3879 = n3878 ? n3877 : n3881;
  /* fppowtf32.vhdl:4400:90  */
  assign n3881 = {1'b0, level0_d1};
  /* fppowtf32.vhdl:4401:23  */
  assign n3883 = {level1_d1, 2'b00};
  /* fppowtf32.vhdl:4401:55  */
  assign n3884 = ps_d1[1]; // extract
  /* fppowtf32.vhdl:4401:45  */
  assign n3885 = n3884 ? n3883 : n3887;
  /* fppowtf32.vhdl:4401:93  */
  assign n3887 = {2'b00, level1_d1};
  /* fppowtf32.vhdl:4402:20  */
  assign n3889 = {level2, 4'b0000};
  /* fppowtf32.vhdl:4402:52  */
  assign n3890 = ps_d1[2]; // extract
  /* fppowtf32.vhdl:4402:42  */
  assign n3891 = n3890 ? n3889 : n3893;
  /* fppowtf32.vhdl:4402:90  */
  assign n3893 = {4'b0000, level2};
  /* fppowtf32.vhdl:4403:20  */
  assign n3895 = {level3, 8'b00000000};
  /* fppowtf32.vhdl:4403:52  */
  assign n3896 = ps_d1[3]; // extract
  /* fppowtf32.vhdl:4403:42  */
  assign n3897 = n3896 ? n3895 : n3899;
  /* fppowtf32.vhdl:4403:90  */
  assign n3899 = {8'b00000000, level3};
  /* fppowtf32.vhdl:4404:20  */
  assign n3901 = {level4, 16'b0000000000000000};
  /* fppowtf32.vhdl:4404:53  */
  assign n3902 = ps_d1[4]; // extract
  /* fppowtf32.vhdl:4404:43  */
  assign n3903 = n3902 ? n3901 : n3905;
  /* fppowtf32.vhdl:4404:92  */
  assign n3905 = {16'b0000000000000000, level4};
  /* fppowtf32.vhdl:4405:15  */
  assign n3906 = level5[40:0]; // extract
  /* fppowtf32.vhdl:4392:10  */
  always @(posedge clk)
    n3907 <= ps;
  /* fppowtf32.vhdl:4392:10  */
  always @(posedge clk)
    n3908 <= level0;
  /* fppowtf32.vhdl:4392:10  */
  always @(posedge clk)
    n3909 <= level1;
endmodule

module intadder_31_freq500_uid69
  (input  clk,
   input  [30:0] x,
   input  [30:0] y,
   input  cin,
   output [30:0] r);
  wire [30:0] rtmp;
  wire [30:0] y_d1;
  wire [30:0] y_d2;
  wire [30:0] y_d3;
  wire [30:0] y_d4;
  wire [30:0] y_d5;
  wire [30:0] y_d6;
  wire [30:0] y_d7;
  wire [30:0] y_d8;
  wire [30:0] y_d9;
  wire [30:0] y_d10;
  wire [30:0] y_d11;
  wire [30:0] y_d12;
  wire [30:0] y_d13;
  wire cin_d1;
  wire cin_d2;
  wire cin_d3;
  wire cin_d4;
  wire cin_d5;
  wire cin_d6;
  wire cin_d7;
  wire cin_d8;
  wire cin_d9;
  wire cin_d10;
  wire cin_d11;
  wire cin_d12;
  wire cin_d13;
  wire [30:0] n3839;
  wire [30:0] n3840;
  wire [30:0] n3841;
  reg [30:0] n3842;
  reg [30:0] n3843;
  reg [30:0] n3844;
  reg [30:0] n3845;
  reg [30:0] n3846;
  reg [30:0] n3847;
  reg [30:0] n3848;
  reg [30:0] n3849;
  reg [30:0] n3850;
  reg [30:0] n3851;
  reg [30:0] n3852;
  reg [30:0] n3853;
  reg [30:0] n3854;
  reg n3855;
  reg n3856;
  reg n3857;
  reg n3858;
  reg n3859;
  reg n3860;
  reg n3861;
  reg n3862;
  reg n3863;
  reg n3864;
  reg n3865;
  reg n3866;
  reg n3867;
  assign r = rtmp; //(module output)
  /* fppowtf32.vhdl:4120:8  */
  assign rtmp = n3841; // (signal)
  /* fppowtf32.vhdl:4122:8  */
  assign y_d1 = n3842; // (signal)
  /* fppowtf32.vhdl:4122:14  */
  assign y_d2 = n3843; // (signal)
  /* fppowtf32.vhdl:4122:20  */
  assign y_d3 = n3844; // (signal)
  /* fppowtf32.vhdl:4122:26  */
  assign y_d4 = n3845; // (signal)
  /* fppowtf32.vhdl:4122:32  */
  assign y_d5 = n3846; // (signal)
  /* fppowtf32.vhdl:4122:38  */
  assign y_d6 = n3847; // (signal)
  /* fppowtf32.vhdl:4122:44  */
  assign y_d7 = n3848; // (signal)
  /* fppowtf32.vhdl:4122:50  */
  assign y_d8 = n3849; // (signal)
  /* fppowtf32.vhdl:4122:56  */
  assign y_d9 = n3850; // (signal)
  /* fppowtf32.vhdl:4122:62  */
  assign y_d10 = n3851; // (signal)
  /* fppowtf32.vhdl:4122:69  */
  assign y_d11 = n3852; // (signal)
  /* fppowtf32.vhdl:4122:76  */
  assign y_d12 = n3853; // (signal)
  /* fppowtf32.vhdl:4122:83  */
  assign y_d13 = n3854; // (signal)
  /* fppowtf32.vhdl:4124:8  */
  assign cin_d1 = n3855; // (signal)
  /* fppowtf32.vhdl:4124:16  */
  assign cin_d2 = n3856; // (signal)
  /* fppowtf32.vhdl:4124:24  */
  assign cin_d3 = n3857; // (signal)
  /* fppowtf32.vhdl:4124:32  */
  assign cin_d4 = n3858; // (signal)
  /* fppowtf32.vhdl:4124:40  */
  assign cin_d5 = n3859; // (signal)
  /* fppowtf32.vhdl:4124:48  */
  assign cin_d6 = n3860; // (signal)
  /* fppowtf32.vhdl:4124:56  */
  assign cin_d7 = n3861; // (signal)
  /* fppowtf32.vhdl:4124:64  */
  assign cin_d8 = n3862; // (signal)
  /* fppowtf32.vhdl:4124:72  */
  assign cin_d9 = n3863; // (signal)
  /* fppowtf32.vhdl:4124:80  */
  assign cin_d10 = n3864; // (signal)
  /* fppowtf32.vhdl:4124:89  */
  assign cin_d11 = n3865; // (signal)
  /* fppowtf32.vhdl:4124:98  */
  assign cin_d12 = n3866; // (signal)
  /* fppowtf32.vhdl:4124:107  */
  assign cin_d13 = n3867; // (signal)
  /* fppowtf32.vhdl:4158:14  */
  assign n3839 = x + y_d13;
  /* fppowtf32.vhdl:4158:22  */
  assign n3840 = {30'b0, cin_d13};  //  uext
  /* fppowtf32.vhdl:4158:22  */
  assign n3841 = n3839 + n3840;
  /* fppowtf32.vhdl:4129:10  */
  always @(posedge clk)
    n3842 <= y;
  /* fppowtf32.vhdl:4129:10  */
  always @(posedge clk)
    n3843 <= y_d1;
  /* fppowtf32.vhdl:4129:10  */
  always @(posedge clk)
    n3844 <= y_d2;
  /* fppowtf32.vhdl:4129:10  */
  always @(posedge clk)
    n3845 <= y_d3;
  /* fppowtf32.vhdl:4129:10  */
  always @(posedge clk)
    n3846 <= y_d4;
  /* fppowtf32.vhdl:4129:10  */
  always @(posedge clk)
    n3847 <= y_d5;
  /* fppowtf32.vhdl:4129:10  */
  always @(posedge clk)
    n3848 <= y_d6;
  /* fppowtf32.vhdl:4129:10  */
  always @(posedge clk)
    n3849 <= y_d7;
  /* fppowtf32.vhdl:4129:10  */
  always @(posedge clk)
    n3850 <= y_d8;
  /* fppowtf32.vhdl:4129:10  */
  always @(posedge clk)
    n3851 <= y_d9;
  /* fppowtf32.vhdl:4129:10  */
  always @(posedge clk)
    n3852 <= y_d10;
  /* fppowtf32.vhdl:4129:10  */
  always @(posedge clk)
    n3853 <= y_d11;
  /* fppowtf32.vhdl:4129:10  */
  always @(posedge clk)
    n3854 <= y_d12;
  /* fppowtf32.vhdl:4129:10  */
  always @(posedge clk)
    n3855 <= cin;
  /* fppowtf32.vhdl:4129:10  */
  always @(posedge clk)
    n3856 <= cin_d1;
  /* fppowtf32.vhdl:4129:10  */
  always @(posedge clk)
    n3857 <= cin_d2;
  /* fppowtf32.vhdl:4129:10  */
  always @(posedge clk)
    n3858 <= cin_d3;
  /* fppowtf32.vhdl:4129:10  */
  always @(posedge clk)
    n3859 <= cin_d4;
  /* fppowtf32.vhdl:4129:10  */
  always @(posedge clk)
    n3860 <= cin_d5;
  /* fppowtf32.vhdl:4129:10  */
  always @(posedge clk)
    n3861 <= cin_d6;
  /* fppowtf32.vhdl:4129:10  */
  always @(posedge clk)
    n3862 <= cin_d7;
  /* fppowtf32.vhdl:4129:10  */
  always @(posedge clk)
    n3863 <= cin_d8;
  /* fppowtf32.vhdl:4129:10  */
  always @(posedge clk)
    n3864 <= cin_d9;
  /* fppowtf32.vhdl:4129:10  */
  always @(posedge clk)
    n3865 <= cin_d10;
  /* fppowtf32.vhdl:4129:10  */
  always @(posedge clk)
    n3866 <= cin_d11;
  /* fppowtf32.vhdl:4129:10  */
  always @(posedge clk)
    n3867 <= cin_d12;
endmodule

module intmultiplier_21x11_24_freq500_uid65
  (input  clk,
   input  [20:0] x,
   input  [10:0] y,
   output [23:0] r);
  wire [20:0] xx;
  wire [10:0] yy;
  wire [10:0] yy_d1;
  wire [10:0] yy_d2;
  wire [10:0] yy_d3;
  wire [10:0] yy_d4;
  wire [10:0] yy_d5;
  wire [10:0] yy_d6;
  wire [10:0] yy_d7;
  wire [10:0] yy_d8;
  wire [10:0] yy_d9;
  wire [10:0] yy_d10;
  wire [10:0] yy_d11;
  wire [31:0] rr;
  wire [31:0] n3793;
  wire [31:0] n3794;
  wire [31:0] n3795;
  wire [23:0] n3796;
  reg [10:0] n3797;
  reg [10:0] n3798;
  reg [10:0] n3799;
  reg [10:0] n3800;
  reg [10:0] n3801;
  reg [10:0] n3802;
  reg [10:0] n3803;
  reg [10:0] n3804;
  reg [10:0] n3805;
  reg [10:0] n3806;
  reg [10:0] n3807;
  assign r = n3796; //(module output)
  /* fppowtf32.vhdl:4059:12  */
  assign yy_d1 = n3797; // (signal)
  /* fppowtf32.vhdl:4059:19  */
  assign yy_d2 = n3798; // (signal)
  /* fppowtf32.vhdl:4059:26  */
  assign yy_d3 = n3799; // (signal)
  /* fppowtf32.vhdl:4059:33  */
  assign yy_d4 = n3800; // (signal)
  /* fppowtf32.vhdl:4059:40  */
  assign yy_d5 = n3801; // (signal)
  /* fppowtf32.vhdl:4059:47  */
  assign yy_d6 = n3802; // (signal)
  /* fppowtf32.vhdl:4059:54  */
  assign yy_d7 = n3803; // (signal)
  /* fppowtf32.vhdl:4059:61  */
  assign yy_d8 = n3804; // (signal)
  /* fppowtf32.vhdl:4059:68  */
  assign yy_d9 = n3805; // (signal)
  /* fppowtf32.vhdl:4059:75  */
  assign yy_d10 = n3806; // (signal)
  /* fppowtf32.vhdl:4059:83  */
  assign yy_d11 = n3807; // (signal)
  /* fppowtf32.vhdl:4061:8  */
  assign rr = n3795; // (signal)
  /* fppowtf32.vhdl:4084:12  */
  assign n3793 = {11'b0, xx};  //  uext
  /* fppowtf32.vhdl:4084:12  */
  assign n3794 = {21'b0, yy_d11};  //  uext
  /* fppowtf32.vhdl:4084:12  */
  assign n3795 = n3793 * n3794; // umul
  /* fppowtf32.vhdl:4085:28  */
  assign n3796 = rr[31:8]; // extract
  /* fppowtf32.vhdl:4066:10  */
  always @(posedge clk)
    n3797 <= yy;
  /* fppowtf32.vhdl:4066:10  */
  always @(posedge clk)
    n3798 <= yy_d1;
  /* fppowtf32.vhdl:4066:10  */
  always @(posedge clk)
    n3799 <= yy_d2;
  /* fppowtf32.vhdl:4066:10  */
  always @(posedge clk)
    n3800 <= yy_d3;
  /* fppowtf32.vhdl:4066:10  */
  always @(posedge clk)
    n3801 <= yy_d4;
  /* fppowtf32.vhdl:4066:10  */
  always @(posedge clk)
    n3802 <= yy_d5;
  /* fppowtf32.vhdl:4066:10  */
  always @(posedge clk)
    n3803 <= yy_d6;
  /* fppowtf32.vhdl:4066:10  */
  always @(posedge clk)
    n3804 <= yy_d7;
  /* fppowtf32.vhdl:4066:10  */
  always @(posedge clk)
    n3805 <= yy_d8;
  /* fppowtf32.vhdl:4066:10  */
  always @(posedge clk)
    n3806 <= yy_d9;
  /* fppowtf32.vhdl:4066:10  */
  always @(posedge clk)
    n3807 <= yy_d10;
endmodule

module intadder_28_freq500_uid60
  (input  clk,
   input  [27:0] x,
   input  [27:0] y,
   input  cin,
   output [27:0] r);
  wire [27:0] rtmp;
  wire cin_d1;
  wire cin_d2;
  wire cin_d3;
  wire cin_d4;
  wire cin_d5;
  wire cin_d6;
  wire cin_d7;
  wire cin_d8;
  wire cin_d9;
  wire cin_d10;
  wire cin_d11;
  wire [27:0] n3763;
  wire [27:0] n3764;
  wire [27:0] n3765;
  reg n3766;
  reg n3767;
  reg n3768;
  reg n3769;
  reg n3770;
  reg n3771;
  reg n3772;
  reg n3773;
  reg n3774;
  reg n3775;
  reg n3776;
  assign r = rtmp; //(module output)
  /* fppowtf32.vhdl:3436:8  */
  assign rtmp = n3765; // (signal)
  /* fppowtf32.vhdl:3438:8  */
  assign cin_d1 = n3766; // (signal)
  /* fppowtf32.vhdl:3438:16  */
  assign cin_d2 = n3767; // (signal)
  /* fppowtf32.vhdl:3438:24  */
  assign cin_d3 = n3768; // (signal)
  /* fppowtf32.vhdl:3438:32  */
  assign cin_d4 = n3769; // (signal)
  /* fppowtf32.vhdl:3438:40  */
  assign cin_d5 = n3770; // (signal)
  /* fppowtf32.vhdl:3438:48  */
  assign cin_d6 = n3771; // (signal)
  /* fppowtf32.vhdl:3438:56  */
  assign cin_d7 = n3772; // (signal)
  /* fppowtf32.vhdl:3438:64  */
  assign cin_d8 = n3773; // (signal)
  /* fppowtf32.vhdl:3438:72  */
  assign cin_d9 = n3774; // (signal)
  /* fppowtf32.vhdl:3438:80  */
  assign cin_d10 = n3775; // (signal)
  /* fppowtf32.vhdl:3438:89  */
  assign cin_d11 = n3776; // (signal)
  /* fppowtf32.vhdl:3457:14  */
  assign n3763 = x + y;
  /* fppowtf32.vhdl:3457:18  */
  assign n3764 = {27'b0, cin_d11};  //  uext
  /* fppowtf32.vhdl:3457:18  */
  assign n3765 = n3763 + n3764;
  /* fppowtf32.vhdl:3443:10  */
  always @(posedge clk)
    n3766 <= cin;
  /* fppowtf32.vhdl:3443:10  */
  always @(posedge clk)
    n3767 <= cin_d1;
  /* fppowtf32.vhdl:3443:10  */
  always @(posedge clk)
    n3768 <= cin_d2;
  /* fppowtf32.vhdl:3443:10  */
  always @(posedge clk)
    n3769 <= cin_d3;
  /* fppowtf32.vhdl:3443:10  */
  always @(posedge clk)
    n3770 <= cin_d4;
  /* fppowtf32.vhdl:3443:10  */
  always @(posedge clk)
    n3771 <= cin_d5;
  /* fppowtf32.vhdl:3443:10  */
  always @(posedge clk)
    n3772 <= cin_d6;
  /* fppowtf32.vhdl:3443:10  */
  always @(posedge clk)
    n3773 <= cin_d7;
  /* fppowtf32.vhdl:3443:10  */
  always @(posedge clk)
    n3774 <= cin_d8;
  /* fppowtf32.vhdl:3443:10  */
  always @(posedge clk)
    n3775 <= cin_d9;
  /* fppowtf32.vhdl:3443:10  */
  always @(posedge clk)
    n3776 <= cin_d10;
endmodule

module intadder_26_freq500_uid57
  (input  clk,
   input  [25:0] x,
   input  [25:0] y,
   input  cin,
   output [25:0] r);
  wire [25:0] rtmp;
  wire [25:0] x_d1;
  wire [25:0] x_d2;
  wire cin_d1;
  wire cin_d2;
  wire cin_d3;
  wire cin_d4;
  wire cin_d5;
  wire cin_d6;
  wire [25:0] n3736;
  wire [25:0] n3737;
  wire [25:0] n3738;
  reg [25:0] n3739;
  reg [25:0] n3740;
  reg n3741;
  reg n3742;
  reg n3743;
  reg n3744;
  reg n3745;
  reg n3746;
  assign r = rtmp; //(module output)
  /* fppowtf32.vhdl:3380:8  */
  assign rtmp = n3738; // (signal)
  /* fppowtf32.vhdl:3382:8  */
  assign x_d1 = n3739; // (signal)
  /* fppowtf32.vhdl:3382:14  */
  assign x_d2 = n3740; // (signal)
  /* fppowtf32.vhdl:3384:8  */
  assign cin_d1 = n3741; // (signal)
  /* fppowtf32.vhdl:3384:16  */
  assign cin_d2 = n3742; // (signal)
  /* fppowtf32.vhdl:3384:24  */
  assign cin_d3 = n3743; // (signal)
  /* fppowtf32.vhdl:3384:32  */
  assign cin_d4 = n3744; // (signal)
  /* fppowtf32.vhdl:3384:40  */
  assign cin_d5 = n3745; // (signal)
  /* fppowtf32.vhdl:3384:48  */
  assign cin_d6 = n3746; // (signal)
  /* fppowtf32.vhdl:3400:17  */
  assign n3736 = x_d2 + y;
  /* fppowtf32.vhdl:3400:21  */
  assign n3737 = {25'b0, cin_d6};  //  uext
  /* fppowtf32.vhdl:3400:21  */
  assign n3738 = n3736 + n3737;
  /* fppowtf32.vhdl:3389:10  */
  always @(posedge clk)
    n3739 <= x;
  /* fppowtf32.vhdl:3389:10  */
  always @(posedge clk)
    n3740 <= x_d1;
  /* fppowtf32.vhdl:3389:10  */
  always @(posedge clk)
    n3741 <= cin;
  /* fppowtf32.vhdl:3389:10  */
  always @(posedge clk)
    n3742 <= cin_d1;
  /* fppowtf32.vhdl:3389:10  */
  always @(posedge clk)
    n3743 <= cin_d2;
  /* fppowtf32.vhdl:3389:10  */
  always @(posedge clk)
    n3744 <= cin_d3;
  /* fppowtf32.vhdl:3389:10  */
  always @(posedge clk)
    n3745 <= cin_d4;
  /* fppowtf32.vhdl:3389:10  */
  always @(posedge clk)
    n3746 <= cin_d5;
endmodule

module rightshifter15_by_max_14_freq500_uid55
  (input  clk,
   input  [14:0] x,
   input  [3:0] s,
   output [28:0] r);
  wire [3:0] ps;
  wire [3:0] ps_d1;
  wire [3:0] ps_d2;
  wire [3:0] ps_d3;
  wire [14:0] level0;
  wire [15:0] level1;
  wire [17:0] level2;
  wire [21:0] level3;
  wire [21:0] level3_d1;
  wire [29:0] level4;
  wire [15:0] n3695;
  wire n3696;
  wire [15:0] n3697;
  wire [15:0] n3699;
  wire [17:0] n3701;
  wire n3702;
  wire [17:0] n3703;
  wire [17:0] n3705;
  wire [21:0] n3707;
  wire n3708;
  wire [21:0] n3709;
  wire [21:0] n3711;
  wire [29:0] n3713;
  wire n3714;
  wire [29:0] n3715;
  wire [29:0] n3717;
  wire [28:0] n3718;
  reg [3:0] n3719;
  reg [3:0] n3720;
  reg [3:0] n3721;
  reg [21:0] n3722;
  assign r = n3718; //(module output)
  /* fppowtf32.vhdl:3317:12  */
  assign ps_d1 = n3719; // (signal)
  /* fppowtf32.vhdl:3317:19  */
  assign ps_d2 = n3720; // (signal)
  /* fppowtf32.vhdl:3317:26  */
  assign ps_d3 = n3721; // (signal)
  /* fppowtf32.vhdl:3321:8  */
  assign level1 = n3697; // (signal)
  /* fppowtf32.vhdl:3323:8  */
  assign level2 = n3703; // (signal)
  /* fppowtf32.vhdl:3325:8  */
  assign level3 = n3709; // (signal)
  /* fppowtf32.vhdl:3325:16  */
  assign level3_d1 = n3722; // (signal)
  /* fppowtf32.vhdl:3327:8  */
  assign level4 = n3715; // (signal)
  /* fppowtf32.vhdl:3341:35  */
  assign n3695 = {1'b0, level0};
  /* fppowtf32.vhdl:3341:54  */
  assign n3696 = ps_d2[0]; // extract
  /* fppowtf32.vhdl:3341:44  */
  assign n3697 = n3696 ? n3695 : n3699;
  /* fppowtf32.vhdl:3341:79  */
  assign n3699 = {level0, 1'b0};
  /* fppowtf32.vhdl:3342:35  */
  assign n3701 = {2'b00, level1};
  /* fppowtf32.vhdl:3342:54  */
  assign n3702 = ps_d2[1]; // extract
  /* fppowtf32.vhdl:3342:44  */
  assign n3703 = n3702 ? n3701 : n3705;
  /* fppowtf32.vhdl:3342:79  */
  assign n3705 = {level1, 2'b00};
  /* fppowtf32.vhdl:3343:35  */
  assign n3707 = {4'b0000, level2};
  /* fppowtf32.vhdl:3343:54  */
  assign n3708 = ps_d2[2]; // extract
  /* fppowtf32.vhdl:3343:44  */
  assign n3709 = n3708 ? n3707 : n3711;
  /* fppowtf32.vhdl:3343:79  */
  assign n3711 = {level2, 4'b0000};
  /* fppowtf32.vhdl:3344:35  */
  assign n3713 = {8'b00000000, level3_d1};
  /* fppowtf32.vhdl:3344:57  */
  assign n3714 = ps_d3[3]; // extract
  /* fppowtf32.vhdl:3344:47  */
  assign n3715 = n3714 ? n3713 : n3717;
  /* fppowtf32.vhdl:3344:85  */
  assign n3717 = {level3_d1, 8'b00000000};
  /* fppowtf32.vhdl:3345:15  */
  assign n3718 = level4[29:1]; // extract
  /* fppowtf32.vhdl:3332:10  */
  always @(posedge clk)
    n3719 <= ps;
  /* fppowtf32.vhdl:3332:10  */
  always @(posedge clk)
    n3720 <= ps_d1;
  /* fppowtf32.vhdl:3332:10  */
  always @(posedge clk)
    n3721 <= ps_d2;
  /* fppowtf32.vhdl:3332:10  */
  always @(posedge clk)
    n3722 <= level3;
endmodule

module normalizer_z_43_35_18_freq500_uid53
  (input  clk,
   input  [42:0] x,
   output [4:0] count,
   output [34:0] r);
  wire [42:0] level5;
  wire count4;
  wire count4_d1;
  wire count4_d2;
  wire [42:0] level4;
  wire [42:0] level4_d1;
  wire count3;
  wire count3_d1;
  wire [41:0] level3;
  wire [41:0] level3_d1;
  wire count2;
  wire count2_d1;
  wire [37:0] level2;
  wire count1;
  wire [35:0] level1;
  wire [35:0] level1_d1;
  wire count0;
  wire count0_d1;
  wire [34:0] level0;
  wire [4:0] scount;
  wire [15:0] n3621;
  wire n3623;
  wire n3624;
  wire n3626;
  wire [42:0] n3627;
  wire [26:0] n3628;
  wire [42:0] n3630;
  wire [7:0] n3632;
  wire n3634;
  wire n3635;
  wire [41:0] n3637;
  wire n3638;
  wire [41:0] n3639;
  wire [34:0] n3640;
  wire [41:0] n3642;
  wire [3:0] n3644;
  wire n3646;
  wire n3647;
  wire [37:0] n3649;
  wire n3650;
  wire [37:0] n3651;
  wire [37:0] n3652;
  wire [1:0] n3654;
  wire n3656;
  wire n3657;
  wire [35:0] n3659;
  wire n3660;
  wire [35:0] n3661;
  wire [35:0] n3662;
  wire n3664;
  wire n3666;
  wire n3667;
  wire [34:0] n3669;
  wire n3670;
  wire [34:0] n3671;
  wire [34:0] n3672;
  wire [1:0] n3673;
  wire [2:0] n3674;
  wire [3:0] n3675;
  wire [4:0] n3676;
  reg n3677;
  reg n3678;
  reg [42:0] n3679;
  reg n3680;
  reg [41:0] n3681;
  reg n3682;
  reg [35:0] n3683;
  reg n3684;
  assign count = scount; //(module output)
  assign r = level0; //(module output)
  /* fppowtf32.vhdl:3229:8  */
  assign count4 = n3624; // (signal)
  /* fppowtf32.vhdl:3229:16  */
  assign count4_d1 = n3677; // (signal)
  /* fppowtf32.vhdl:3229:27  */
  assign count4_d2 = n3678; // (signal)
  /* fppowtf32.vhdl:3231:8  */
  assign level4 = n3627; // (signal)
  /* fppowtf32.vhdl:3231:16  */
  assign level4_d1 = n3679; // (signal)
  /* fppowtf32.vhdl:3233:8  */
  assign count3 = n3635; // (signal)
  /* fppowtf32.vhdl:3233:16  */
  assign count3_d1 = n3680; // (signal)
  /* fppowtf32.vhdl:3235:8  */
  assign level3 = n3639; // (signal)
  /* fppowtf32.vhdl:3235:16  */
  assign level3_d1 = n3681; // (signal)
  /* fppowtf32.vhdl:3237:8  */
  assign count2 = n3647; // (signal)
  /* fppowtf32.vhdl:3237:16  */
  assign count2_d1 = n3682; // (signal)
  /* fppowtf32.vhdl:3239:8  */
  assign level2 = n3651; // (signal)
  /* fppowtf32.vhdl:3241:8  */
  assign count1 = n3657; // (signal)
  /* fppowtf32.vhdl:3243:8  */
  assign level1 = n3661; // (signal)
  /* fppowtf32.vhdl:3243:16  */
  assign level1_d1 = n3683; // (signal)
  /* fppowtf32.vhdl:3245:8  */
  assign count0 = n3667; // (signal)
  /* fppowtf32.vhdl:3245:16  */
  assign count0_d1 = n3684; // (signal)
  /* fppowtf32.vhdl:3247:8  */
  assign level0 = n3671; // (signal)
  /* fppowtf32.vhdl:3249:8  */
  assign scount = n3676; // (signal)
  /* fppowtf32.vhdl:3266:28  */
  assign n3621 = level5[42:27]; // extract
  /* fppowtf32.vhdl:3266:43  */
  assign n3623 = n3621 == 16'b0000000000000000;
  /* fppowtf32.vhdl:3266:17  */
  assign n3624 = n3623 ? 1'b1 : 1'b0;
  /* fppowtf32.vhdl:3267:44  */
  assign n3626 = ~count4;
  /* fppowtf32.vhdl:3267:33  */
  assign n3627 = n3626 ? level5 : n3630;
  /* fppowtf32.vhdl:3267:60  */
  assign n3628 = level5[26:0]; // extract
  /* fppowtf32.vhdl:3267:74  */
  assign n3630 = {n3628, 16'b0000000000000000};
  /* fppowtf32.vhdl:3269:31  */
  assign n3632 = level4_d1[42:35]; // extract
  /* fppowtf32.vhdl:3269:46  */
  assign n3634 = n3632 == 8'b00000000;
  /* fppowtf32.vhdl:3269:17  */
  assign n3635 = n3634 ? 1'b1 : 1'b0;
  /* fppowtf32.vhdl:3270:22  */
  assign n3637 = level4_d1[42:1]; // extract
  /* fppowtf32.vhdl:3270:47  */
  assign n3638 = ~count3;
  /* fppowtf32.vhdl:3270:36  */
  assign n3639 = n3638 ? n3637 : n3642;
  /* fppowtf32.vhdl:3270:66  */
  assign n3640 = level4_d1[34:0]; // extract
  /* fppowtf32.vhdl:3270:80  */
  assign n3642 = {n3640, 7'b0000000};
  /* fppowtf32.vhdl:3272:28  */
  assign n3644 = level3[41:38]; // extract
  /* fppowtf32.vhdl:3272:43  */
  assign n3646 = n3644 == 4'b0000;
  /* fppowtf32.vhdl:3272:17  */
  assign n3647 = n3646 ? 1'b1 : 1'b0;
  /* fppowtf32.vhdl:3273:22  */
  assign n3649 = level3_d1[41:4]; // extract
  /* fppowtf32.vhdl:3273:50  */
  assign n3650 = ~count2_d1;
  /* fppowtf32.vhdl:3273:36  */
  assign n3651 = n3650 ? n3649 : n3652;
  /* fppowtf32.vhdl:3273:69  */
  assign n3652 = level3_d1[37:0]; // extract
  /* fppowtf32.vhdl:3275:28  */
  assign n3654 = level2[37:36]; // extract
  /* fppowtf32.vhdl:3275:43  */
  assign n3656 = n3654 == 2'b00;
  /* fppowtf32.vhdl:3275:17  */
  assign n3657 = n3656 ? 1'b1 : 1'b0;
  /* fppowtf32.vhdl:3276:19  */
  assign n3659 = level2[37:2]; // extract
  /* fppowtf32.vhdl:3276:44  */
  assign n3660 = ~count1;
  /* fppowtf32.vhdl:3276:33  */
  assign n3661 = n3660 ? n3659 : n3662;
  /* fppowtf32.vhdl:3276:60  */
  assign n3662 = level2[35:0]; // extract
  /* fppowtf32.vhdl:3278:28  */
  assign n3664 = level1[35]; // extract
  /* fppowtf32.vhdl:3278:43  */
  assign n3666 = n3664 == 1'b0;
  /* fppowtf32.vhdl:3278:17  */
  assign n3667 = n3666 ? 1'b1 : 1'b0;
  /* fppowtf32.vhdl:3279:22  */
  assign n3669 = level1_d1[35:1]; // extract
  /* fppowtf32.vhdl:3279:50  */
  assign n3670 = ~count0_d1;
  /* fppowtf32.vhdl:3279:36  */
  assign n3671 = n3670 ? n3669 : n3672;
  /* fppowtf32.vhdl:3279:69  */
  assign n3672 = level1_d1[34:0]; // extract
  /* fppowtf32.vhdl:3282:24  */
  assign n3673 = {count4_d2, count3_d1};
  /* fppowtf32.vhdl:3282:36  */
  assign n3674 = {n3673, count2_d1};
  /* fppowtf32.vhdl:3282:48  */
  assign n3675 = {n3674, count1};
  /* fppowtf32.vhdl:3282:57  */
  assign n3676 = {n3675, count0};
  /* fppowtf32.vhdl:3254:10  */
  always @(posedge clk)
    n3677 <= count4;
  /* fppowtf32.vhdl:3254:10  */
  always @(posedge clk)
    n3678 <= count4_d1;
  /* fppowtf32.vhdl:3254:10  */
  always @(posedge clk)
    n3679 <= level4;
  /* fppowtf32.vhdl:3254:10  */
  always @(posedge clk)
    n3680 <= count3;
  /* fppowtf32.vhdl:3254:10  */
  always @(posedge clk)
    n3681 <= level3;
  /* fppowtf32.vhdl:3254:10  */
  always @(posedge clk)
    n3682 <= count2;
  /* fppowtf32.vhdl:3254:10  */
  always @(posedge clk)
    n3683 <= level1;
  /* fppowtf32.vhdl:3254:10  */
  always @(posedge clk)
    n3684 <= count0;
endmodule

module intadder_43_freq500_uid51
  (input  clk,
   input  [42:0] x,
   input  [42:0] y,
   input  cin,
   output [42:0] r);
  wire cin_0;
  wire cin_0_d1;
  wire cin_0_d2;
  wire cin_0_d3;
  wire cin_0_d4;
  wire cin_0_d5;
  wire cin_0_d6;
  wire cin_0_d7;
  wire [25:0] x_0;
  wire [25:0] x_0_d1;
  wire [25:0] x_0_d2;
  wire [25:0] x_0_d3;
  wire [25:0] x_0_d4;
  wire [25:0] x_0_d5;
  wire [25:0] x_0_d6;
  wire [25:0] y_0;
  wire [25:0] y_0_d1;
  wire [25:0] s_0;
  wire [24:0] r_0;
  wire [24:0] r_0_d1;
  wire cin_1;
  wire cin_1_d1;
  wire [18:0] x_1;
  wire [18:0] x_1_d1;
  wire [18:0] x_1_d2;
  wire [18:0] x_1_d3;
  wire [18:0] x_1_d4;
  wire [18:0] x_1_d5;
  wire [18:0] x_1_d6;
  wire [18:0] x_1_d7;
  wire [18:0] y_1;
  wire [18:0] y_1_d1;
  wire [18:0] y_1_d2;
  wire [18:0] s_1;
  wire [17:0] r_1;
  wire [24:0] n3559;
  wire [25:0] n3561;
  wire [24:0] n3562;
  wire [25:0] n3564;
  wire [25:0] n3565;
  wire [25:0] n3566;
  wire [25:0] n3567;
  wire [24:0] n3568;
  wire n3569;
  wire [17:0] n3570;
  wire [18:0] n3572;
  wire [17:0] n3573;
  wire [18:0] n3575;
  wire [18:0] n3576;
  wire [18:0] n3577;
  wire [18:0] n3578;
  wire [17:0] n3579;
  wire [42:0] n3580;
  reg n3581;
  reg n3582;
  reg n3583;
  reg n3584;
  reg n3585;
  reg n3586;
  reg n3587;
  reg [25:0] n3588;
  reg [25:0] n3589;
  reg [25:0] n3590;
  reg [25:0] n3591;
  reg [25:0] n3592;
  reg [25:0] n3593;
  reg [25:0] n3594;
  reg [24:0] n3595;
  reg n3596;
  reg [18:0] n3597;
  reg [18:0] n3598;
  reg [18:0] n3599;
  reg [18:0] n3600;
  reg [18:0] n3601;
  reg [18:0] n3602;
  reg [18:0] n3603;
  reg [18:0] n3604;
  reg [18:0] n3605;
  assign r = n3580; //(module output)
  /* fppowtf32.vhdl:3132:15  */
  assign cin_0_d1 = n3581; // (signal)
  /* fppowtf32.vhdl:3132:25  */
  assign cin_0_d2 = n3582; // (signal)
  /* fppowtf32.vhdl:3132:35  */
  assign cin_0_d3 = n3583; // (signal)
  /* fppowtf32.vhdl:3132:45  */
  assign cin_0_d4 = n3584; // (signal)
  /* fppowtf32.vhdl:3132:55  */
  assign cin_0_d5 = n3585; // (signal)
  /* fppowtf32.vhdl:3132:65  */
  assign cin_0_d6 = n3586; // (signal)
  /* fppowtf32.vhdl:3132:75  */
  assign cin_0_d7 = n3587; // (signal)
  /* fppowtf32.vhdl:3134:8  */
  assign x_0 = n3561; // (signal)
  /* fppowtf32.vhdl:3134:13  */
  assign x_0_d1 = n3588; // (signal)
  /* fppowtf32.vhdl:3134:21  */
  assign x_0_d2 = n3589; // (signal)
  /* fppowtf32.vhdl:3134:29  */
  assign x_0_d3 = n3590; // (signal)
  /* fppowtf32.vhdl:3134:37  */
  assign x_0_d4 = n3591; // (signal)
  /* fppowtf32.vhdl:3134:45  */
  assign x_0_d5 = n3592; // (signal)
  /* fppowtf32.vhdl:3134:53  */
  assign x_0_d6 = n3593; // (signal)
  /* fppowtf32.vhdl:3136:8  */
  assign y_0 = n3564; // (signal)
  /* fppowtf32.vhdl:3136:13  */
  assign y_0_d1 = n3594; // (signal)
  /* fppowtf32.vhdl:3138:8  */
  assign s_0 = n3567; // (signal)
  /* fppowtf32.vhdl:3140:8  */
  assign r_0 = n3568; // (signal)
  /* fppowtf32.vhdl:3140:13  */
  assign r_0_d1 = n3595; // (signal)
  /* fppowtf32.vhdl:3142:8  */
  assign cin_1 = n3569; // (signal)
  /* fppowtf32.vhdl:3142:15  */
  assign cin_1_d1 = n3596; // (signal)
  /* fppowtf32.vhdl:3144:8  */
  assign x_1 = n3572; // (signal)
  /* fppowtf32.vhdl:3144:13  */
  assign x_1_d1 = n3597; // (signal)
  /* fppowtf32.vhdl:3144:21  */
  assign x_1_d2 = n3598; // (signal)
  /* fppowtf32.vhdl:3144:29  */
  assign x_1_d3 = n3599; // (signal)
  /* fppowtf32.vhdl:3144:37  */
  assign x_1_d4 = n3600; // (signal)
  /* fppowtf32.vhdl:3144:45  */
  assign x_1_d5 = n3601; // (signal)
  /* fppowtf32.vhdl:3144:53  */
  assign x_1_d6 = n3602; // (signal)
  /* fppowtf32.vhdl:3144:61  */
  assign x_1_d7 = n3603; // (signal)
  /* fppowtf32.vhdl:3146:8  */
  assign y_1 = n3575; // (signal)
  /* fppowtf32.vhdl:3146:13  */
  assign y_1_d1 = n3604; // (signal)
  /* fppowtf32.vhdl:3146:21  */
  assign y_1_d2 = n3605; // (signal)
  /* fppowtf32.vhdl:3148:8  */
  assign s_1 = n3578; // (signal)
  /* fppowtf32.vhdl:3150:8  */
  assign r_1 = n3579; // (signal)
  /* fppowtf32.vhdl:3184:18  */
  assign n3559 = x[24:0]; // extract
  /* fppowtf32.vhdl:3184:15  */
  assign n3561 = {1'b0, n3559};
  /* fppowtf32.vhdl:3185:18  */
  assign n3562 = y[24:0]; // extract
  /* fppowtf32.vhdl:3185:15  */
  assign n3564 = {1'b0, n3562};
  /* fppowtf32.vhdl:3186:18  */
  assign n3565 = x_0_d6 + y_0_d1;
  /* fppowtf32.vhdl:3186:27  */
  assign n3566 = {25'b0, cin_0_d7};  //  uext
  /* fppowtf32.vhdl:3186:27  */
  assign n3567 = n3565 + n3566;
  /* fppowtf32.vhdl:3187:14  */
  assign n3568 = s_0[24:0]; // extract
  /* fppowtf32.vhdl:3188:16  */
  assign n3569 = s_0[25]; // extract
  /* fppowtf32.vhdl:3189:18  */
  assign n3570 = x[42:25]; // extract
  /* fppowtf32.vhdl:3189:15  */
  assign n3572 = {1'b0, n3570};
  /* fppowtf32.vhdl:3190:18  */
  assign n3573 = y[42:25]; // extract
  /* fppowtf32.vhdl:3190:15  */
  assign n3575 = {1'b0, n3573};
  /* fppowtf32.vhdl:3191:18  */
  assign n3576 = x_1_d7 + y_1_d2;
  /* fppowtf32.vhdl:3191:27  */
  assign n3577 = {18'b0, cin_1_d1};  //  uext
  /* fppowtf32.vhdl:3191:27  */
  assign n3578 = n3576 + n3577;
  /* fppowtf32.vhdl:3192:14  */
  assign n3579 = s_1[17:0]; // extract
  /* fppowtf32.vhdl:3193:13  */
  assign n3580 = {r_1, r_0_d1};
  /* fppowtf32.vhdl:3155:10  */
  always @(posedge clk)
    n3581 <= cin_0;
  /* fppowtf32.vhdl:3155:10  */
  always @(posedge clk)
    n3582 <= cin_0_d1;
  /* fppowtf32.vhdl:3155:10  */
  always @(posedge clk)
    n3583 <= cin_0_d2;
  /* fppowtf32.vhdl:3155:10  */
  always @(posedge clk)
    n3584 <= cin_0_d3;
  /* fppowtf32.vhdl:3155:10  */
  always @(posedge clk)
    n3585 <= cin_0_d4;
  /* fppowtf32.vhdl:3155:10  */
  always @(posedge clk)
    n3586 <= cin_0_d5;
  /* fppowtf32.vhdl:3155:10  */
  always @(posedge clk)
    n3587 <= cin_0_d6;
  /* fppowtf32.vhdl:3155:10  */
  always @(posedge clk)
    n3588 <= x_0;
  /* fppowtf32.vhdl:3155:10  */
  always @(posedge clk)
    n3589 <= x_0_d1;
  /* fppowtf32.vhdl:3155:10  */
  always @(posedge clk)
    n3590 <= x_0_d2;
  /* fppowtf32.vhdl:3155:10  */
  always @(posedge clk)
    n3591 <= x_0_d3;
  /* fppowtf32.vhdl:3155:10  */
  always @(posedge clk)
    n3592 <= x_0_d4;
  /* fppowtf32.vhdl:3155:10  */
  always @(posedge clk)
    n3593 <= x_0_d5;
  /* fppowtf32.vhdl:3155:10  */
  always @(posedge clk)
    n3594 <= y_0;
  /* fppowtf32.vhdl:3155:10  */
  always @(posedge clk)
    n3595 <= r_0;
  /* fppowtf32.vhdl:3155:10  */
  always @(posedge clk)
    n3596 <= cin_1;
  /* fppowtf32.vhdl:3155:10  */
  always @(posedge clk)
    n3597 <= x_1;
  /* fppowtf32.vhdl:3155:10  */
  always @(posedge clk)
    n3598 <= x_1_d1;
  /* fppowtf32.vhdl:3155:10  */
  always @(posedge clk)
    n3599 <= x_1_d2;
  /* fppowtf32.vhdl:3155:10  */
  always @(posedge clk)
    n3600 <= x_1_d3;
  /* fppowtf32.vhdl:3155:10  */
  always @(posedge clk)
    n3601 <= x_1_d4;
  /* fppowtf32.vhdl:3155:10  */
  always @(posedge clk)
    n3602 <= x_1_d5;
  /* fppowtf32.vhdl:3155:10  */
  always @(posedge clk)
    n3603 <= x_1_d6;
  /* fppowtf32.vhdl:3155:10  */
  always @(posedge clk)
    n3604 <= y_1;
  /* fppowtf32.vhdl:3155:10  */
  always @(posedge clk)
    n3605 <= y_1_d1;
endmodule

module fixrealkcm_freq500_uid39
  (input  clk,
   input  [7:0] x,
   output [31:0] r);
  wire [4:0] fixrealkcm_freq500_uid39_a0;
  wire [31:0] fixrealkcm_freq500_uid39_t0;
  wire [31:0] fixrealkcm_freq500_uid39_t0_copy43;
  wire [31:0] fixrealkcm_freq500_uid39_t0_copy43_d1;
  wire bh40_w0_0;
  wire bh40_w1_0;
  wire bh40_w2_0;
  wire bh40_w3_0;
  wire bh40_w4_0;
  wire bh40_w5_0;
  wire bh40_w6_0;
  wire bh40_w7_0;
  wire bh40_w8_0;
  wire bh40_w9_0;
  wire bh40_w10_0;
  wire bh40_w11_0;
  wire bh40_w12_0;
  wire bh40_w13_0;
  wire bh40_w14_0;
  wire bh40_w15_0;
  wire bh40_w16_0;
  wire bh40_w17_0;
  wire bh40_w18_0;
  wire bh40_w19_0;
  wire bh40_w20_0;
  wire bh40_w21_0;
  wire bh40_w22_0;
  wire bh40_w23_0;
  wire bh40_w24_0;
  wire bh40_w25_0;
  wire bh40_w26_0;
  wire bh40_w27_0;
  wire bh40_w28_0;
  wire bh40_w29_0;
  wire bh40_w30_0;
  wire bh40_w31_0;
  wire [2:0] fixrealkcm_freq500_uid39_a1;
  wire [26:0] fixrealkcm_freq500_uid39_t1;
  wire [26:0] fixrealkcm_freq500_uid39_t1_copy46;
  wire [26:0] fixrealkcm_freq500_uid39_t1_copy46_d1;
  wire bh40_w0_1;
  wire bh40_w1_1;
  wire bh40_w2_1;
  wire bh40_w3_1;
  wire bh40_w4_1;
  wire bh40_w5_1;
  wire bh40_w6_1;
  wire bh40_w7_1;
  wire bh40_w8_1;
  wire bh40_w9_1;
  wire bh40_w10_1;
  wire bh40_w11_1;
  wire bh40_w12_1;
  wire bh40_w13_1;
  wire bh40_w14_1;
  wire bh40_w15_1;
  wire bh40_w16_1;
  wire bh40_w17_1;
  wire bh40_w18_1;
  wire bh40_w19_1;
  wire bh40_w20_1;
  wire bh40_w21_1;
  wire bh40_w22_1;
  wire bh40_w23_1;
  wire bh40_w24_1;
  wire bh40_w25_1;
  wire bh40_w26_1;
  wire [31:0] bitheapfinaladd_bh40_in0;
  wire [31:0] bitheapfinaladd_bh40_in1;
  wire bitheapfinaladd_bh40_cin;
  wire [31:0] bitheapfinaladd_bh40_out;
  wire [31:0] bitheapresult_bh40;
  wire [31:0] outres;
  wire [4:0] n3396;
  wire [31:0] fixrealkcm_freq500_uid39_table0_n3397;
  wire n3400;
  wire n3401;
  wire n3402;
  wire n3403;
  wire n3404;
  wire n3405;
  wire n3406;
  wire n3407;
  wire n3408;
  wire n3409;
  wire n3410;
  wire n3411;
  wire n3412;
  wire n3413;
  wire n3414;
  wire n3415;
  wire n3416;
  wire n3417;
  wire n3418;
  wire n3419;
  wire n3420;
  wire n3421;
  wire n3422;
  wire n3423;
  wire n3424;
  wire n3425;
  wire n3426;
  wire n3427;
  wire n3428;
  wire n3429;
  wire n3430;
  wire n3431;
  wire [2:0] n3432;
  wire [26:0] fixrealkcm_freq500_uid39_table1_n3433;
  wire n3436;
  wire n3437;
  wire n3438;
  wire n3439;
  wire n3440;
  wire n3441;
  wire n3442;
  wire n3443;
  wire n3444;
  wire n3445;
  wire n3446;
  wire n3447;
  wire n3448;
  wire n3449;
  wire n3450;
  wire n3451;
  wire n3452;
  wire n3453;
  wire n3454;
  wire n3455;
  wire n3456;
  wire n3457;
  wire n3458;
  wire n3459;
  wire n3460;
  wire n3461;
  wire n3462;
  wire [1:0] n3464;
  wire [2:0] n3465;
  wire [3:0] n3466;
  wire [4:0] n3467;
  wire [5:0] n3468;
  wire [6:0] n3469;
  wire [7:0] n3470;
  wire [8:0] n3471;
  wire [9:0] n3472;
  wire [10:0] n3473;
  wire [11:0] n3474;
  wire [12:0] n3475;
  wire [13:0] n3476;
  wire [14:0] n3477;
  wire [15:0] n3478;
  wire [16:0] n3479;
  wire [17:0] n3480;
  wire [18:0] n3481;
  wire [19:0] n3482;
  wire [20:0] n3483;
  wire [21:0] n3484;
  wire [22:0] n3485;
  wire [23:0] n3486;
  wire [24:0] n3487;
  wire [25:0] n3488;
  wire [26:0] n3489;
  wire [27:0] n3490;
  wire [28:0] n3491;
  wire [29:0] n3492;
  wire [30:0] n3493;
  wire [31:0] n3494;
  wire [5:0] n3496;
  wire [6:0] n3497;
  wire [7:0] n3498;
  wire [8:0] n3499;
  wire [9:0] n3500;
  wire [10:0] n3501;
  wire [11:0] n3502;
  wire [12:0] n3503;
  wire [13:0] n3504;
  wire [14:0] n3505;
  wire [15:0] n3506;
  wire [16:0] n3507;
  wire [17:0] n3508;
  wire [18:0] n3509;
  wire [19:0] n3510;
  wire [20:0] n3511;
  wire [21:0] n3512;
  wire [22:0] n3513;
  wire [23:0] n3514;
  wire [24:0] n3515;
  wire [25:0] n3516;
  wire [26:0] n3517;
  wire [27:0] n3518;
  wire [28:0] n3519;
  wire [29:0] n3520;
  wire [30:0] n3521;
  wire [31:0] n3522;
  wire [31:0] bitheapfinaladd_bh40_n3524;
  reg [31:0] n3527;
  reg [26:0] n3528;
  assign r = outres; //(module output)
  /* fppowtf32.vhdl:2860:8  */
  assign fixrealkcm_freq500_uid39_a0 = n3396; // (signal)
  /* fppowtf32.vhdl:2862:8  */
  assign fixrealkcm_freq500_uid39_t0 = fixrealkcm_freq500_uid39_t0_copy43_d1; // (signal)
  /* fppowtf32.vhdl:2864:8  */
  assign fixrealkcm_freq500_uid39_t0_copy43 = fixrealkcm_freq500_uid39_table0_n3397; // (signal)
  /* fppowtf32.vhdl:2864:44  */
  assign fixrealkcm_freq500_uid39_t0_copy43_d1 = n3527; // (signal)
  /* fppowtf32.vhdl:2866:8  */
  assign bh40_w0_0 = n3400; // (signal)
  /* fppowtf32.vhdl:2868:8  */
  assign bh40_w1_0 = n3401; // (signal)
  /* fppowtf32.vhdl:2870:8  */
  assign bh40_w2_0 = n3402; // (signal)
  /* fppowtf32.vhdl:2872:8  */
  assign bh40_w3_0 = n3403; // (signal)
  /* fppowtf32.vhdl:2874:8  */
  assign bh40_w4_0 = n3404; // (signal)
  /* fppowtf32.vhdl:2876:8  */
  assign bh40_w5_0 = n3405; // (signal)
  /* fppowtf32.vhdl:2878:8  */
  assign bh40_w6_0 = n3406; // (signal)
  /* fppowtf32.vhdl:2880:8  */
  assign bh40_w7_0 = n3407; // (signal)
  /* fppowtf32.vhdl:2882:8  */
  assign bh40_w8_0 = n3408; // (signal)
  /* fppowtf32.vhdl:2884:8  */
  assign bh40_w9_0 = n3409; // (signal)
  /* fppowtf32.vhdl:2886:8  */
  assign bh40_w10_0 = n3410; // (signal)
  /* fppowtf32.vhdl:2888:8  */
  assign bh40_w11_0 = n3411; // (signal)
  /* fppowtf32.vhdl:2890:8  */
  assign bh40_w12_0 = n3412; // (signal)
  /* fppowtf32.vhdl:2892:8  */
  assign bh40_w13_0 = n3413; // (signal)
  /* fppowtf32.vhdl:2894:8  */
  assign bh40_w14_0 = n3414; // (signal)
  /* fppowtf32.vhdl:2896:8  */
  assign bh40_w15_0 = n3415; // (signal)
  /* fppowtf32.vhdl:2898:8  */
  assign bh40_w16_0 = n3416; // (signal)
  /* fppowtf32.vhdl:2900:8  */
  assign bh40_w17_0 = n3417; // (signal)
  /* fppowtf32.vhdl:2902:8  */
  assign bh40_w18_0 = n3418; // (signal)
  /* fppowtf32.vhdl:2904:8  */
  assign bh40_w19_0 = n3419; // (signal)
  /* fppowtf32.vhdl:2906:8  */
  assign bh40_w20_0 = n3420; // (signal)
  /* fppowtf32.vhdl:2908:8  */
  assign bh40_w21_0 = n3421; // (signal)
  /* fppowtf32.vhdl:2910:8  */
  assign bh40_w22_0 = n3422; // (signal)
  /* fppowtf32.vhdl:2912:8  */
  assign bh40_w23_0 = n3423; // (signal)
  /* fppowtf32.vhdl:2914:8  */
  assign bh40_w24_0 = n3424; // (signal)
  /* fppowtf32.vhdl:2916:8  */
  assign bh40_w25_0 = n3425; // (signal)
  /* fppowtf32.vhdl:2918:8  */
  assign bh40_w26_0 = n3426; // (signal)
  /* fppowtf32.vhdl:2920:8  */
  assign bh40_w27_0 = n3427; // (signal)
  /* fppowtf32.vhdl:2922:8  */
  assign bh40_w28_0 = n3428; // (signal)
  /* fppowtf32.vhdl:2924:8  */
  assign bh40_w29_0 = n3429; // (signal)
  /* fppowtf32.vhdl:2926:8  */
  assign bh40_w30_0 = n3430; // (signal)
  /* fppowtf32.vhdl:3085:35  */
  assign bh40_w31_0 = n3431; // (signal)
  /* fppowtf32.vhdl:2930:8  */
  assign fixrealkcm_freq500_uid39_a1 = n3432; // (signal)
  /* fppowtf32.vhdl:2932:8  */
  assign fixrealkcm_freq500_uid39_t1 = fixrealkcm_freq500_uid39_t1_copy46_d1; // (signal)
  /* fppowtf32.vhdl:2934:8  */
  assign fixrealkcm_freq500_uid39_t1_copy46 = fixrealkcm_freq500_uid39_table1_n3433; // (signal)
  /* fppowtf32.vhdl:2934:44  */
  assign fixrealkcm_freq500_uid39_t1_copy46_d1 = n3528; // (signal)
  /* fppowtf32.vhdl:2936:8  */
  assign bh40_w0_1 = n3436; // (signal)
  /* fppowtf32.vhdl:2938:8  */
  assign bh40_w1_1 = n3437; // (signal)
  /* fppowtf32.vhdl:2940:8  */
  assign bh40_w2_1 = n3438; // (signal)
  /* fppowtf32.vhdl:2942:8  */
  assign bh40_w3_1 = n3439; // (signal)
  /* fppowtf32.vhdl:2944:8  */
  assign bh40_w4_1 = n3440; // (signal)
  /* fppowtf32.vhdl:2946:8  */
  assign bh40_w5_1 = n3441; // (signal)
  /* fppowtf32.vhdl:2948:8  */
  assign bh40_w6_1 = n3442; // (signal)
  /* fppowtf32.vhdl:2950:8  */
  assign bh40_w7_1 = n3443; // (signal)
  /* fppowtf32.vhdl:2952:8  */
  assign bh40_w8_1 = n3444; // (signal)
  /* fppowtf32.vhdl:2954:8  */
  assign bh40_w9_1 = n3445; // (signal)
  /* fppowtf32.vhdl:2956:8  */
  assign bh40_w10_1 = n3446; // (signal)
  /* fppowtf32.vhdl:2958:8  */
  assign bh40_w11_1 = n3447; // (signal)
  /* fppowtf32.vhdl:2960:8  */
  assign bh40_w12_1 = n3448; // (signal)
  /* fppowtf32.vhdl:2962:8  */
  assign bh40_w13_1 = n3449; // (signal)
  /* fppowtf32.vhdl:2964:8  */
  assign bh40_w14_1 = n3450; // (signal)
  /* fppowtf32.vhdl:2966:8  */
  assign bh40_w15_1 = n3451; // (signal)
  /* fppowtf32.vhdl:2968:8  */
  assign bh40_w16_1 = n3452; // (signal)
  /* fppowtf32.vhdl:2970:8  */
  assign bh40_w17_1 = n3453; // (signal)
  /* fppowtf32.vhdl:2972:8  */
  assign bh40_w18_1 = n3454; // (signal)
  /* fppowtf32.vhdl:2974:8  */
  assign bh40_w19_1 = n3455; // (signal)
  /* fppowtf32.vhdl:2976:8  */
  assign bh40_w20_1 = n3456; // (signal)
  /* fppowtf32.vhdl:2978:8  */
  assign bh40_w21_1 = n3457; // (signal)
  /* fppowtf32.vhdl:2980:8  */
  assign bh40_w22_1 = n3458; // (signal)
  /* fppowtf32.vhdl:2982:8  */
  assign bh40_w23_1 = n3459; // (signal)
  /* fppowtf32.vhdl:2984:8  */
  assign bh40_w24_1 = n3460; // (signal)
  /* fppowtf32.vhdl:2986:8  */
  assign bh40_w25_1 = n3461; // (signal)
  /* fppowtf32.vhdl:2988:8  */
  assign bh40_w26_1 = n3462; // (signal)
  /* fppowtf32.vhdl:2990:8  */
  assign bitheapfinaladd_bh40_in0 = n3494; // (signal)
  /* fppowtf32.vhdl:2992:8  */
  assign bitheapfinaladd_bh40_in1 = n3522; // (signal)
  /* fppowtf32.vhdl:2994:8  */
  assign bitheapfinaladd_bh40_cin = 1'b0; // (signal)
  /* fppowtf32.vhdl:2996:8  */
  assign bitheapfinaladd_bh40_out = bitheapfinaladd_bh40_n3524; // (signal)
  /* fppowtf32.vhdl:2998:8  */
  assign bitheapresult_bh40 = bitheapfinaladd_bh40_out; // (signal)
  /* fppowtf32.vhdl:3000:8  */
  assign outres = bitheapresult_bh40; // (signal)
  /* fppowtf32.vhdl:3011:36  */
  assign n3396 = x[7:3]; // extract
  /* fppowtf32.vhdl:3012:4  */
  fixrealkcm_freq500_uid39_t0_freq500_uid42 fixrealkcm_freq500_uid39_table0 (
    .x(fixrealkcm_freq500_uid39_a0),
    .y(fixrealkcm_freq500_uid39_table0_n3397));
  /* fppowtf32.vhdl:3016:44  */
  assign n3400 = fixrealkcm_freq500_uid39_t0[0]; // extract
  /* fppowtf32.vhdl:3017:44  */
  assign n3401 = fixrealkcm_freq500_uid39_t0[1]; // extract
  /* fppowtf32.vhdl:3018:44  */
  assign n3402 = fixrealkcm_freq500_uid39_t0[2]; // extract
  /* fppowtf32.vhdl:3019:44  */
  assign n3403 = fixrealkcm_freq500_uid39_t0[3]; // extract
  /* fppowtf32.vhdl:3020:44  */
  assign n3404 = fixrealkcm_freq500_uid39_t0[4]; // extract
  /* fppowtf32.vhdl:3021:44  */
  assign n3405 = fixrealkcm_freq500_uid39_t0[5]; // extract
  /* fppowtf32.vhdl:3022:44  */
  assign n3406 = fixrealkcm_freq500_uid39_t0[6]; // extract
  /* fppowtf32.vhdl:3023:44  */
  assign n3407 = fixrealkcm_freq500_uid39_t0[7]; // extract
  /* fppowtf32.vhdl:3024:44  */
  assign n3408 = fixrealkcm_freq500_uid39_t0[8]; // extract
  /* fppowtf32.vhdl:3025:44  */
  assign n3409 = fixrealkcm_freq500_uid39_t0[9]; // extract
  /* fppowtf32.vhdl:3026:45  */
  assign n3410 = fixrealkcm_freq500_uid39_t0[10]; // extract
  /* fppowtf32.vhdl:3027:45  */
  assign n3411 = fixrealkcm_freq500_uid39_t0[11]; // extract
  /* fppowtf32.vhdl:3028:45  */
  assign n3412 = fixrealkcm_freq500_uid39_t0[12]; // extract
  /* fppowtf32.vhdl:3029:45  */
  assign n3413 = fixrealkcm_freq500_uid39_t0[13]; // extract
  /* fppowtf32.vhdl:3030:45  */
  assign n3414 = fixrealkcm_freq500_uid39_t0[14]; // extract
  /* fppowtf32.vhdl:3031:45  */
  assign n3415 = fixrealkcm_freq500_uid39_t0[15]; // extract
  /* fppowtf32.vhdl:3032:45  */
  assign n3416 = fixrealkcm_freq500_uid39_t0[16]; // extract
  /* fppowtf32.vhdl:3033:45  */
  assign n3417 = fixrealkcm_freq500_uid39_t0[17]; // extract
  /* fppowtf32.vhdl:3034:45  */
  assign n3418 = fixrealkcm_freq500_uid39_t0[18]; // extract
  /* fppowtf32.vhdl:3035:45  */
  assign n3419 = fixrealkcm_freq500_uid39_t0[19]; // extract
  /* fppowtf32.vhdl:3036:45  */
  assign n3420 = fixrealkcm_freq500_uid39_t0[20]; // extract
  /* fppowtf32.vhdl:3037:45  */
  assign n3421 = fixrealkcm_freq500_uid39_t0[21]; // extract
  /* fppowtf32.vhdl:3038:45  */
  assign n3422 = fixrealkcm_freq500_uid39_t0[22]; // extract
  /* fppowtf32.vhdl:3039:45  */
  assign n3423 = fixrealkcm_freq500_uid39_t0[23]; // extract
  /* fppowtf32.vhdl:3040:45  */
  assign n3424 = fixrealkcm_freq500_uid39_t0[24]; // extract
  /* fppowtf32.vhdl:3041:45  */
  assign n3425 = fixrealkcm_freq500_uid39_t0[25]; // extract
  /* fppowtf32.vhdl:3042:45  */
  assign n3426 = fixrealkcm_freq500_uid39_t0[26]; // extract
  /* fppowtf32.vhdl:3043:45  */
  assign n3427 = fixrealkcm_freq500_uid39_t0[27]; // extract
  /* fppowtf32.vhdl:3044:45  */
  assign n3428 = fixrealkcm_freq500_uid39_t0[28]; // extract
  /* fppowtf32.vhdl:3045:45  */
  assign n3429 = fixrealkcm_freq500_uid39_t0[29]; // extract
  /* fppowtf32.vhdl:3046:45  */
  assign n3430 = fixrealkcm_freq500_uid39_t0[30]; // extract
  /* fppowtf32.vhdl:3047:45  */
  assign n3431 = fixrealkcm_freq500_uid39_t0[31]; // extract
  /* fppowtf32.vhdl:3048:36  */
  assign n3432 = x[2:0]; // extract
  /* fppowtf32.vhdl:3049:4  */
  fixrealkcm_freq500_uid39_t1_freq500_uid45 fixrealkcm_freq500_uid39_table1 (
    .x(fixrealkcm_freq500_uid39_a1),
    .y(fixrealkcm_freq500_uid39_table1_n3433));
  /* fppowtf32.vhdl:3053:44  */
  assign n3436 = fixrealkcm_freq500_uid39_t1[0]; // extract
  /* fppowtf32.vhdl:3054:44  */
  assign n3437 = fixrealkcm_freq500_uid39_t1[1]; // extract
  /* fppowtf32.vhdl:3055:44  */
  assign n3438 = fixrealkcm_freq500_uid39_t1[2]; // extract
  /* fppowtf32.vhdl:3056:44  */
  assign n3439 = fixrealkcm_freq500_uid39_t1[3]; // extract
  /* fppowtf32.vhdl:3057:44  */
  assign n3440 = fixrealkcm_freq500_uid39_t1[4]; // extract
  /* fppowtf32.vhdl:3058:44  */
  assign n3441 = fixrealkcm_freq500_uid39_t1[5]; // extract
  /* fppowtf32.vhdl:3059:44  */
  assign n3442 = fixrealkcm_freq500_uid39_t1[6]; // extract
  /* fppowtf32.vhdl:3060:44  */
  assign n3443 = fixrealkcm_freq500_uid39_t1[7]; // extract
  /* fppowtf32.vhdl:3061:44  */
  assign n3444 = fixrealkcm_freq500_uid39_t1[8]; // extract
  /* fppowtf32.vhdl:3062:44  */
  assign n3445 = fixrealkcm_freq500_uid39_t1[9]; // extract
  /* fppowtf32.vhdl:3063:45  */
  assign n3446 = fixrealkcm_freq500_uid39_t1[10]; // extract
  /* fppowtf32.vhdl:3064:45  */
  assign n3447 = fixrealkcm_freq500_uid39_t1[11]; // extract
  /* fppowtf32.vhdl:3065:45  */
  assign n3448 = fixrealkcm_freq500_uid39_t1[12]; // extract
  /* fppowtf32.vhdl:3066:45  */
  assign n3449 = fixrealkcm_freq500_uid39_t1[13]; // extract
  /* fppowtf32.vhdl:3067:45  */
  assign n3450 = fixrealkcm_freq500_uid39_t1[14]; // extract
  /* fppowtf32.vhdl:3068:45  */
  assign n3451 = fixrealkcm_freq500_uid39_t1[15]; // extract
  /* fppowtf32.vhdl:3069:45  */
  assign n3452 = fixrealkcm_freq500_uid39_t1[16]; // extract
  /* fppowtf32.vhdl:3070:45  */
  assign n3453 = fixrealkcm_freq500_uid39_t1[17]; // extract
  /* fppowtf32.vhdl:3071:45  */
  assign n3454 = fixrealkcm_freq500_uid39_t1[18]; // extract
  /* fppowtf32.vhdl:3072:45  */
  assign n3455 = fixrealkcm_freq500_uid39_t1[19]; // extract
  /* fppowtf32.vhdl:3073:45  */
  assign n3456 = fixrealkcm_freq500_uid39_t1[20]; // extract
  /* fppowtf32.vhdl:3074:45  */
  assign n3457 = fixrealkcm_freq500_uid39_t1[21]; // extract
  /* fppowtf32.vhdl:3075:45  */
  assign n3458 = fixrealkcm_freq500_uid39_t1[22]; // extract
  /* fppowtf32.vhdl:3076:45  */
  assign n3459 = fixrealkcm_freq500_uid39_t1[23]; // extract
  /* fppowtf32.vhdl:3077:45  */
  assign n3460 = fixrealkcm_freq500_uid39_t1[24]; // extract
  /* fppowtf32.vhdl:3078:45  */
  assign n3461 = fixrealkcm_freq500_uid39_t1[25]; // extract
  /* fppowtf32.vhdl:3079:45  */
  assign n3462 = fixrealkcm_freq500_uid39_t1[26]; // extract
  /* fppowtf32.vhdl:3085:48  */
  assign n3464 = {bh40_w31_0, bh40_w30_0};
  /* fppowtf32.vhdl:3085:61  */
  assign n3465 = {n3464, bh40_w29_0};
  /* fppowtf32.vhdl:3085:74  */
  assign n3466 = {n3465, bh40_w28_0};
  /* fppowtf32.vhdl:3085:87  */
  assign n3467 = {n3466, bh40_w27_0};
  /* fppowtf32.vhdl:3085:100  */
  assign n3468 = {n3467, bh40_w26_1};
  /* fppowtf32.vhdl:3085:113  */
  assign n3469 = {n3468, bh40_w25_1};
  /* fppowtf32.vhdl:3085:126  */
  assign n3470 = {n3469, bh40_w24_1};
  /* fppowtf32.vhdl:3085:139  */
  assign n3471 = {n3470, bh40_w23_1};
  /* fppowtf32.vhdl:3085:152  */
  assign n3472 = {n3471, bh40_w22_1};
  /* fppowtf32.vhdl:3085:165  */
  assign n3473 = {n3472, bh40_w21_1};
  /* fppowtf32.vhdl:3085:178  */
  assign n3474 = {n3473, bh40_w20_1};
  /* fppowtf32.vhdl:3085:191  */
  assign n3475 = {n3474, bh40_w19_1};
  /* fppowtf32.vhdl:3085:204  */
  assign n3476 = {n3475, bh40_w18_1};
  /* fppowtf32.vhdl:3085:217  */
  assign n3477 = {n3476, bh40_w17_1};
  /* fppowtf32.vhdl:3085:230  */
  assign n3478 = {n3477, bh40_w16_1};
  /* fppowtf32.vhdl:3085:243  */
  assign n3479 = {n3478, bh40_w15_1};
  /* fppowtf32.vhdl:3085:256  */
  assign n3480 = {n3479, bh40_w14_1};
  /* fppowtf32.vhdl:3085:269  */
  assign n3481 = {n3480, bh40_w13_1};
  /* fppowtf32.vhdl:3085:282  */
  assign n3482 = {n3481, bh40_w12_1};
  /* fppowtf32.vhdl:3085:295  */
  assign n3483 = {n3482, bh40_w11_1};
  /* fppowtf32.vhdl:3085:308  */
  assign n3484 = {n3483, bh40_w10_1};
  /* fppowtf32.vhdl:3085:321  */
  assign n3485 = {n3484, bh40_w9_1};
  /* fppowtf32.vhdl:3085:333  */
  assign n3486 = {n3485, bh40_w8_1};
  /* fppowtf32.vhdl:3085:345  */
  assign n3487 = {n3486, bh40_w7_1};
  /* fppowtf32.vhdl:3085:357  */
  assign n3488 = {n3487, bh40_w6_1};
  /* fppowtf32.vhdl:3085:369  */
  assign n3489 = {n3488, bh40_w5_1};
  /* fppowtf32.vhdl:3085:381  */
  assign n3490 = {n3489, bh40_w4_1};
  /* fppowtf32.vhdl:3085:393  */
  assign n3491 = {n3490, bh40_w3_1};
  /* fppowtf32.vhdl:3085:405  */
  assign n3492 = {n3491, bh40_w2_1};
  /* fppowtf32.vhdl:3085:417  */
  assign n3493 = {n3492, bh40_w1_1};
  /* fppowtf32.vhdl:3085:429  */
  assign n3494 = {n3493, bh40_w0_1};
  /* fppowtf32.vhdl:3086:60  */
  assign n3496 = {5'b00000, bh40_w26_0};
  /* fppowtf32.vhdl:3086:73  */
  assign n3497 = {n3496, bh40_w25_0};
  /* fppowtf32.vhdl:3086:86  */
  assign n3498 = {n3497, bh40_w24_0};
  /* fppowtf32.vhdl:3086:99  */
  assign n3499 = {n3498, bh40_w23_0};
  /* fppowtf32.vhdl:3086:112  */
  assign n3500 = {n3499, bh40_w22_0};
  /* fppowtf32.vhdl:3086:125  */
  assign n3501 = {n3500, bh40_w21_0};
  /* fppowtf32.vhdl:3086:138  */
  assign n3502 = {n3501, bh40_w20_0};
  /* fppowtf32.vhdl:3086:151  */
  assign n3503 = {n3502, bh40_w19_0};
  /* fppowtf32.vhdl:3086:164  */
  assign n3504 = {n3503, bh40_w18_0};
  /* fppowtf32.vhdl:3086:177  */
  assign n3505 = {n3504, bh40_w17_0};
  /* fppowtf32.vhdl:3086:190  */
  assign n3506 = {n3505, bh40_w16_0};
  /* fppowtf32.vhdl:3086:203  */
  assign n3507 = {n3506, bh40_w15_0};
  /* fppowtf32.vhdl:3086:216  */
  assign n3508 = {n3507, bh40_w14_0};
  /* fppowtf32.vhdl:3086:229  */
  assign n3509 = {n3508, bh40_w13_0};
  /* fppowtf32.vhdl:3086:242  */
  assign n3510 = {n3509, bh40_w12_0};
  /* fppowtf32.vhdl:3086:255  */
  assign n3511 = {n3510, bh40_w11_0};
  /* fppowtf32.vhdl:3086:268  */
  assign n3512 = {n3511, bh40_w10_0};
  /* fppowtf32.vhdl:3086:281  */
  assign n3513 = {n3512, bh40_w9_0};
  /* fppowtf32.vhdl:3086:293  */
  assign n3514 = {n3513, bh40_w8_0};
  /* fppowtf32.vhdl:3086:305  */
  assign n3515 = {n3514, bh40_w7_0};
  /* fppowtf32.vhdl:3086:317  */
  assign n3516 = {n3515, bh40_w6_0};
  /* fppowtf32.vhdl:3086:329  */
  assign n3517 = {n3516, bh40_w5_0};
  /* fppowtf32.vhdl:3086:341  */
  assign n3518 = {n3517, bh40_w4_0};
  /* fppowtf32.vhdl:3086:353  */
  assign n3519 = {n3518, bh40_w3_0};
  /* fppowtf32.vhdl:3086:365  */
  assign n3520 = {n3519, bh40_w2_0};
  /* fppowtf32.vhdl:3086:377  */
  assign n3521 = {n3520, bh40_w1_0};
  /* fppowtf32.vhdl:3086:389  */
  assign n3522 = {n3521, bh40_w0_0};
  /* fppowtf32.vhdl:3089:4  */
  intadder_32_freq500_uid49 bitheapfinaladd_bh40 (
    .clk(clk),
    .x(bitheapfinaladd_bh40_in0),
    .y(bitheapfinaladd_bh40_in1),
    .cin(bitheapfinaladd_bh40_cin),
    .r(bitheapfinaladd_bh40_n3524));
  /* fppowtf32.vhdl:3005:10  */
  always @(posedge clk)
    n3527 <= fixrealkcm_freq500_uid39_t0_copy43;
  /* fppowtf32.vhdl:3005:10  */
  always @(posedge clk)
    n3528 <= fixrealkcm_freq500_uid39_t1_copy46;
endmodule

module intadder_35_freq500_uid37
  (input  clk,
   input  [34:0] x,
   input  [34:0] y,
   input  cin,
   output [34:0] r);
  wire [34:0] rtmp;
  wire [34:0] x_d1;
  wire [34:0] x_d2;
  wire [34:0] x_d3;
  wire [34:0] x_d4;
  wire cin_d1;
  wire cin_d2;
  wire cin_d3;
  wire cin_d4;
  wire cin_d5;
  wire cin_d6;
  wire [34:0] n3376;
  wire [34:0] n3377;
  wire [34:0] n3378;
  reg [34:0] n3379;
  reg [34:0] n3380;
  reg [34:0] n3381;
  reg [34:0] n3382;
  reg n3383;
  reg n3384;
  reg n3385;
  reg n3386;
  reg n3387;
  reg n3388;
  assign r = rtmp; //(module output)
  /* fppowtf32.vhdl:2739:8  */
  assign rtmp = n3378; // (signal)
  /* fppowtf32.vhdl:2741:8  */
  assign x_d1 = n3379; // (signal)
  /* fppowtf32.vhdl:2741:14  */
  assign x_d2 = n3380; // (signal)
  /* fppowtf32.vhdl:2741:20  */
  assign x_d3 = n3381; // (signal)
  /* fppowtf32.vhdl:2741:26  */
  assign x_d4 = n3382; // (signal)
  /* fppowtf32.vhdl:2743:8  */
  assign cin_d1 = n3383; // (signal)
  /* fppowtf32.vhdl:2743:16  */
  assign cin_d2 = n3384; // (signal)
  /* fppowtf32.vhdl:2743:24  */
  assign cin_d3 = n3385; // (signal)
  /* fppowtf32.vhdl:2743:32  */
  assign cin_d4 = n3386; // (signal)
  /* fppowtf32.vhdl:2743:40  */
  assign cin_d5 = n3387; // (signal)
  /* fppowtf32.vhdl:2743:48  */
  assign cin_d6 = n3388; // (signal)
  /* fppowtf32.vhdl:2761:17  */
  assign n3376 = x_d4 + y;
  /* fppowtf32.vhdl:2761:21  */
  assign n3377 = {34'b0, cin_d6};  //  uext
  /* fppowtf32.vhdl:2761:21  */
  assign n3378 = n3376 + n3377;
  /* fppowtf32.vhdl:2748:10  */
  always @(posedge clk)
    n3379 <= x;
  /* fppowtf32.vhdl:2748:10  */
  always @(posedge clk)
    n3380 <= x_d1;
  /* fppowtf32.vhdl:2748:10  */
  always @(posedge clk)
    n3381 <= x_d2;
  /* fppowtf32.vhdl:2748:10  */
  always @(posedge clk)
    n3382 <= x_d3;
  /* fppowtf32.vhdl:2748:10  */
  always @(posedge clk)
    n3383 <= cin;
  /* fppowtf32.vhdl:2748:10  */
  always @(posedge clk)
    n3384 <= cin_d1;
  /* fppowtf32.vhdl:2748:10  */
  always @(posedge clk)
    n3385 <= cin_d2;
  /* fppowtf32.vhdl:2748:10  */
  always @(posedge clk)
    n3386 <= cin_d3;
  /* fppowtf32.vhdl:2748:10  */
  always @(posedge clk)
    n3387 <= cin_d4;
  /* fppowtf32.vhdl:2748:10  */
  always @(posedge clk)
    n3388 <= cin_d5;
endmodule

module intadder_35_freq500_uid34
  (input  clk,
   input  [34:0] x,
   input  [34:0] y,
   input  cin,
   output [34:0] r);
  wire cin_1;
  wire cin_1_d1;
  wire cin_1_d2;
  wire [35:0] x_1;
  wire [35:0] x_1_d1;
  wire [35:0] x_1_d2;
  wire [35:0] y_1;
  wire [35:0] y_1_d1;
  wire [35:0] s_1;
  wire [34:0] r_1;
  wire [35:0] n3349;
  wire [35:0] n3351;
  wire [35:0] n3352;
  wire [35:0] n3353;
  wire [35:0] n3354;
  wire [34:0] n3355;
  reg n3356;
  reg n3357;
  reg [35:0] n3358;
  reg [35:0] n3359;
  reg [35:0] n3360;
  assign r = r_1; //(module output)
  /* fppowtf32.vhdl:2678:15  */
  assign cin_1_d1 = n3356; // (signal)
  /* fppowtf32.vhdl:2678:25  */
  assign cin_1_d2 = n3357; // (signal)
  /* fppowtf32.vhdl:2680:8  */
  assign x_1 = n3349; // (signal)
  /* fppowtf32.vhdl:2680:13  */
  assign x_1_d1 = n3358; // (signal)
  /* fppowtf32.vhdl:2680:21  */
  assign x_1_d2 = n3359; // (signal)
  /* fppowtf32.vhdl:2682:8  */
  assign y_1 = n3351; // (signal)
  /* fppowtf32.vhdl:2682:13  */
  assign y_1_d1 = n3360; // (signal)
  /* fppowtf32.vhdl:2684:8  */
  assign s_1 = n3354; // (signal)
  /* fppowtf32.vhdl:2686:8  */
  assign r_1 = n3355; // (signal)
  /* fppowtf32.vhdl:2700:15  */
  assign n3349 = {1'b0, x};
  /* fppowtf32.vhdl:2701:15  */
  assign n3351 = {1'b0, y};
  /* fppowtf32.vhdl:2702:18  */
  assign n3352 = x_1_d2 + y_1_d1;
  /* fppowtf32.vhdl:2702:27  */
  assign n3353 = {35'b0, cin_1_d2};  //  uext
  /* fppowtf32.vhdl:2702:27  */
  assign n3354 = n3352 + n3353;
  /* fppowtf32.vhdl:2703:14  */
  assign n3355 = s_1[34:0]; // extract
  /* fppowtf32.vhdl:2691:10  */
  always @(posedge clk)
    n3356 <= cin_1;
  /* fppowtf32.vhdl:2691:10  */
  always @(posedge clk)
    n3357 <= cin_1_d1;
  /* fppowtf32.vhdl:2691:10  */
  always @(posedge clk)
    n3358 <= x_1;
  /* fppowtf32.vhdl:2691:10  */
  always @(posedge clk)
    n3359 <= x_1_d1;
  /* fppowtf32.vhdl:2691:10  */
  always @(posedge clk)
    n3360 <= y_1;
endmodule

module logtable1_freq500_uid30
  (input  [5:0] x,
   output [28:0] y);
  wire [28:0] y0;
  wire [28:0] y1;
  wire n3145;
  wire n3148;
  wire n3151;
  wire n3154;
  wire n3157;
  wire n3160;
  wire n3163;
  wire n3166;
  wire n3169;
  wire n3172;
  wire n3175;
  wire n3178;
  wire n3181;
  wire n3184;
  wire n3187;
  wire n3190;
  wire n3193;
  wire n3196;
  wire n3199;
  wire n3202;
  wire n3205;
  wire n3208;
  wire n3211;
  wire n3214;
  wire n3217;
  wire n3220;
  wire n3223;
  wire n3226;
  wire n3229;
  wire n3232;
  wire n3235;
  wire n3238;
  wire n3241;
  wire n3244;
  wire n3247;
  wire n3250;
  wire n3253;
  wire n3256;
  wire n3259;
  wire n3262;
  wire n3265;
  wire n3268;
  wire n3271;
  wire n3274;
  wire n3277;
  wire n3280;
  wire n3283;
  wire n3286;
  wire n3289;
  wire n3292;
  wire n3295;
  wire n3298;
  wire n3301;
  wire n3304;
  wire n3307;
  wire n3310;
  wire n3313;
  wire n3316;
  wire n3319;
  wire n3322;
  wire n3325;
  wire n3328;
  wire n3331;
  wire n3334;
  wire [63:0] n3336;
  reg [28:0] n3337;
  assign y = y1; //(module output)
  /* fppowtf32.vhdl:622:8  */
  assign y0 = n3337; // (signal)
  /* fppowtf32.vhdl:624:8  */
  assign y1 = y0; // (signal)
  /* fppowtf32.vhdl:628:39  */
  assign n3145 = x == 6'b000000;
  /* fppowtf32.vhdl:629:39  */
  assign n3148 = x == 6'b000001;
  /* fppowtf32.vhdl:630:39  */
  assign n3151 = x == 6'b000010;
  /* fppowtf32.vhdl:631:39  */
  assign n3154 = x == 6'b000011;
  /* fppowtf32.vhdl:632:39  */
  assign n3157 = x == 6'b000100;
  /* fppowtf32.vhdl:633:39  */
  assign n3160 = x == 6'b000101;
  /* fppowtf32.vhdl:634:39  */
  assign n3163 = x == 6'b000110;
  /* fppowtf32.vhdl:635:39  */
  assign n3166 = x == 6'b000111;
  /* fppowtf32.vhdl:636:39  */
  assign n3169 = x == 6'b001000;
  /* fppowtf32.vhdl:637:39  */
  assign n3172 = x == 6'b001001;
  /* fppowtf32.vhdl:638:39  */
  assign n3175 = x == 6'b001010;
  /* fppowtf32.vhdl:639:39  */
  assign n3178 = x == 6'b001011;
  /* fppowtf32.vhdl:640:39  */
  assign n3181 = x == 6'b001100;
  /* fppowtf32.vhdl:641:39  */
  assign n3184 = x == 6'b001101;
  /* fppowtf32.vhdl:642:39  */
  assign n3187 = x == 6'b001110;
  /* fppowtf32.vhdl:643:39  */
  assign n3190 = x == 6'b001111;
  /* fppowtf32.vhdl:644:39  */
  assign n3193 = x == 6'b010000;
  /* fppowtf32.vhdl:645:39  */
  assign n3196 = x == 6'b010001;
  /* fppowtf32.vhdl:646:39  */
  assign n3199 = x == 6'b010010;
  /* fppowtf32.vhdl:647:39  */
  assign n3202 = x == 6'b010011;
  /* fppowtf32.vhdl:648:39  */
  assign n3205 = x == 6'b010100;
  /* fppowtf32.vhdl:649:39  */
  assign n3208 = x == 6'b010101;
  /* fppowtf32.vhdl:650:39  */
  assign n3211 = x == 6'b010110;
  /* fppowtf32.vhdl:651:39  */
  assign n3214 = x == 6'b010111;
  /* fppowtf32.vhdl:652:39  */
  assign n3217 = x == 6'b011000;
  /* fppowtf32.vhdl:653:39  */
  assign n3220 = x == 6'b011001;
  /* fppowtf32.vhdl:654:39  */
  assign n3223 = x == 6'b011010;
  /* fppowtf32.vhdl:655:39  */
  assign n3226 = x == 6'b011011;
  /* fppowtf32.vhdl:656:39  */
  assign n3229 = x == 6'b011100;
  /* fppowtf32.vhdl:657:39  */
  assign n3232 = x == 6'b011101;
  /* fppowtf32.vhdl:658:39  */
  assign n3235 = x == 6'b011110;
  /* fppowtf32.vhdl:659:39  */
  assign n3238 = x == 6'b011111;
  /* fppowtf32.vhdl:660:39  */
  assign n3241 = x == 6'b100000;
  /* fppowtf32.vhdl:661:39  */
  assign n3244 = x == 6'b100001;
  /* fppowtf32.vhdl:662:39  */
  assign n3247 = x == 6'b100010;
  /* fppowtf32.vhdl:663:39  */
  assign n3250 = x == 6'b100011;
  /* fppowtf32.vhdl:664:39  */
  assign n3253 = x == 6'b100100;
  /* fppowtf32.vhdl:665:39  */
  assign n3256 = x == 6'b100101;
  /* fppowtf32.vhdl:666:39  */
  assign n3259 = x == 6'b100110;
  /* fppowtf32.vhdl:667:39  */
  assign n3262 = x == 6'b100111;
  /* fppowtf32.vhdl:668:39  */
  assign n3265 = x == 6'b101000;
  /* fppowtf32.vhdl:669:39  */
  assign n3268 = x == 6'b101001;
  /* fppowtf32.vhdl:670:39  */
  assign n3271 = x == 6'b101010;
  /* fppowtf32.vhdl:671:39  */
  assign n3274 = x == 6'b101011;
  /* fppowtf32.vhdl:672:39  */
  assign n3277 = x == 6'b101100;
  /* fppowtf32.vhdl:673:39  */
  assign n3280 = x == 6'b101101;
  /* fppowtf32.vhdl:674:39  */
  assign n3283 = x == 6'b101110;
  /* fppowtf32.vhdl:675:39  */
  assign n3286 = x == 6'b101111;
  /* fppowtf32.vhdl:676:39  */
  assign n3289 = x == 6'b110000;
  /* fppowtf32.vhdl:677:39  */
  assign n3292 = x == 6'b110001;
  /* fppowtf32.vhdl:678:39  */
  assign n3295 = x == 6'b110010;
  /* fppowtf32.vhdl:679:39  */
  assign n3298 = x == 6'b110011;
  /* fppowtf32.vhdl:680:39  */
  assign n3301 = x == 6'b110100;
  /* fppowtf32.vhdl:681:39  */
  assign n3304 = x == 6'b110101;
  /* fppowtf32.vhdl:682:39  */
  assign n3307 = x == 6'b110110;
  /* fppowtf32.vhdl:683:39  */
  assign n3310 = x == 6'b110111;
  /* fppowtf32.vhdl:684:39  */
  assign n3313 = x == 6'b111000;
  /* fppowtf32.vhdl:685:39  */
  assign n3316 = x == 6'b111001;
  /* fppowtf32.vhdl:686:39  */
  assign n3319 = x == 6'b111010;
  /* fppowtf32.vhdl:687:39  */
  assign n3322 = x == 6'b111011;
  /* fppowtf32.vhdl:688:39  */
  assign n3325 = x == 6'b111100;
  /* fppowtf32.vhdl:689:39  */
  assign n3328 = x == 6'b111101;
  /* fppowtf32.vhdl:690:39  */
  assign n3331 = x == 6'b111110;
  /* fppowtf32.vhdl:691:39  */
  assign n3334 = x == 6'b111111;
  assign n3336 = {n3334, n3331, n3328, n3325, n3322, n3319, n3316, n3313, n3310, n3307, n3304, n3301, n3298, n3295, n3292, n3289, n3286, n3283, n3280, n3277, n3274, n3271, n3268, n3265, n3262, n3259, n3256, n3253, n3250, n3247, n3244, n3241, n3238, n3235, n3232, n3229, n3226, n3223, n3220, n3217, n3214, n3211, n3208, n3205, n3202, n3199, n3196, n3193, n3190, n3187, n3184, n3181, n3178, n3175, n3172, n3169, n3166, n3163, n3160, n3157, n3154, n3151, n3148, n3145};
  /* fppowtf32.vhdl:627:4  */
  always @*
    case (n3336)
      64'b1000000000000000000000000000000000000000000000000000000000000000: n3337 = 29'b11111101111001010110011110010;
      64'b0100000000000000000000000000000000000000000000000000000000000000: n3337 = 29'b11111001110101011100101110010;
      64'b0010000000000000000000000000000000000000000000000000000000000000: n3337 = 29'b11110101110001100111000110000;
      64'b0001000000000000000000000000000000000000000000000000000000000000: n3337 = 29'b11110001101101110101100101100;
      64'b0000100000000000000000000000000000000000000000000000000000000000: n3337 = 29'b11101101101010001000001100100;
      64'b0000010000000000000000000000000000000000000000000000000000000000: n3337 = 29'b11101001100110011110111010111;
      64'b0000001000000000000000000000000000000000000000000000000000000000: n3337 = 29'b11100101100010111001110000101;
      64'b0000000100000000000000000000000000000000000000000000000000000000: n3337 = 29'b11100001011111011000101101011;
      64'b0000000010000000000000000000000000000000000000000000000000000000: n3337 = 29'b11011101011011111011110001010;
      64'b0000000001000000000000000000000000000000000000000000000000000000: n3337 = 29'b11011001011000100010111100000;
      64'b0000000000100000000000000000000000000000000000000000000000000000: n3337 = 29'b11010101010101001110001101100;
      64'b0000000000010000000000000000000000000000000000000000000000000000: n3337 = 29'b11010001010001111101100101101;
      64'b0000000000001000000000000000000000000000000000000000000000000000: n3337 = 29'b11001101001110110001000100010;
      64'b0000000000000100000000000000000000000000000000000000000000000000: n3337 = 29'b11001001001011101000101001010;
      64'b0000000000000010000000000000000000000000000000000000000000000000: n3337 = 29'b11000101001000100100010100100;
      64'b0000000000000001000000000000000000000000000000000000000000000000: n3337 = 29'b11000001000101100100000101110;
      64'b0000000000000000100000000000000000000000000000000000000000000000: n3337 = 29'b10111101000010100111111101001;
      64'b0000000000000000010000000000000000000000000000000000000000000000: n3337 = 29'b10111000111111101111111010010;
      64'b0000000000000000001000000000000000000000000000000000000000000000: n3337 = 29'b10110100111100111011111101001;
      64'b0000000000000000000100000000000000000000000000000000000000000000: n3337 = 29'b10110000111010001100000101100;
      64'b0000000000000000000010000000000000000000000000000000000000000000: n3337 = 29'b10101100110111100000010011100;
      64'b0000000000000000000001000000000000000000000000000000000000000000: n3337 = 29'b10101000110100111000100110110;
      64'b0000000000000000000000100000000000000000000000000000000000000000: n3337 = 29'b10100100110010010100111111001;
      64'b0000000000000000000000010000000000000000000000000000000000000000: n3337 = 29'b10100000101111110101011100110;
      64'b0000000000000000000000001000000000000000000000000000000000000000: n3337 = 29'b10011100101101011001111111001;
      64'b0000000000000000000000000100000000000000000000000000000000000000: n3337 = 29'b10011000101011000010100110100;
      64'b0000000000000000000000000010000000000000000000000000000000000000: n3337 = 29'b10010100101000101111010010100;
      64'b0000000000000000000000000001000000000000000000000000000000000000: n3337 = 29'b10010000100110100000000011000;
      64'b0000000000000000000000000000100000000000000000000000000000000000: n3337 = 29'b10001100100100010100111000000;
      64'b0000000000000000000000000000010000000000000000000000000000000000: n3337 = 29'b10001000100010001101110001010;
      64'b0000000000000000000000000000001000000000000000000000000000000000: n3337 = 29'b10000100100000001010101110110;
      64'b0000000000000000000000000000000100000000000000000000000000000000: n3337 = 29'b10000000011110001011110000010;
      64'b0000000000000000000000000000000010000000000000000000000000000000: n3337 = 29'b01111110011101001101110010100;
      64'b0000000000000000000000000000000001000000000000000000000000000000: n3337 = 29'b01111010011011010100111001110;
      64'b0000000000000000000000000000000000100000000000000000000000000000: n3337 = 29'b01110110011001100000000100110;
      64'b0000000000000000000000000000000000010000000000000000000000000000: n3337 = 29'b01110010010111101111010011100;
      64'b0000000000000000000000000000000000001000000000000000000000000000: n3337 = 29'b01101110010110000010100101100;
      64'b0000000000000000000000000000000000000100000000000000000000000000: n3337 = 29'b01101010010100011001111011000;
      64'b0000000000000000000000000000000000000010000000000000000000000000: n3337 = 29'b01100110010010110101010011110;
      64'b0000000000000000000000000000000000000001000000000000000000000000: n3337 = 29'b01100010010001010100101111100;
      64'b0000000000000000000000000000000000000000100000000000000000000000: n3337 = 29'b01011110001111111000001110010;
      64'b0000000000000000000000000000000000000000010000000000000000000000: n3337 = 29'b01011010001110011111101111111;
      64'b0000000000000000000000000000000000000000001000000000000000000000: n3337 = 29'b01010110001101001011010100010;
      64'b0000000000000000000000000000000000000000000100000000000000000000: n3337 = 29'b01010010001011111010111011000;
      64'b0000000000000000000000000000000000000000000010000000000000000000: n3337 = 29'b01001110001010101110100100011;
      64'b0000000000000000000000000000000000000000000001000000000000000000: n3337 = 29'b01001010001001100110010000000;
      64'b0000000000000000000000000000000000000000000000100000000000000000: n3337 = 29'b01000110001000100001111101111;
      64'b0000000000000000000000000000000000000000000000010000000000000000: n3337 = 29'b01000010000111100001101101110;
      64'b0000000000000000000000000000000000000000000000001000000000000000: n3337 = 29'b00111110000110100101011111110;
      64'b0000000000000000000000000000000000000000000000000100000000000000: n3337 = 29'b00111010000101101101010011011;
      64'b0000000000000000000000000000000000000000000000000010000000000000: n3337 = 29'b00110110000100111001001000110;
      64'b0000000000000000000000000000000000000000000000000001000000000000: n3337 = 29'b00110010000100001000111111110;
      64'b0000000000000000000000000000000000000000000000000000100000000000: n3337 = 29'b00101110000011011100111000001;
      64'b0000000000000000000000000000000000000000000000000000010000000000: n3337 = 29'b00101010000010110100110001111;
      64'b0000000000000000000000000000000000000000000000000000001000000000: n3337 = 29'b00100110000010010000101100110;
      64'b0000000000000000000000000000000000000000000000000000000100000000: n3337 = 29'b00100010000001110000101000110;
      64'b0000000000000000000000000000000000000000000000000000000010000000: n3337 = 29'b00011110000001010100100101110;
      64'b0000000000000000000000000000000000000000000000000000000001000000: n3337 = 29'b00011010000000111100100011100;
      64'b0000000000000000000000000000000000000000000000000000000000100000: n3337 = 29'b00010110000000101000100001111;
      64'b0000000000000000000000000000000000000000000000000000000000010000: n3337 = 29'b00010010000000011000100000111;
      64'b0000000000000000000000000000000000000000000000000000000000001000: n3337 = 29'b00001110000000001100100000011;
      64'b0000000000000000000000000000000000000000000000000000000000000100: n3337 = 29'b00001010000000000100100000001;
      64'b0000000000000000000000000000000000000000000000000000000000000010: n3337 = 29'b00000110000000000000100000000;
      64'b0000000000000000000000000000000000000000000000000000000000000001: n3337 = 29'b00000010000000000000100000000;
      default: n3337 = 29'bX;
    endcase
endmodule

module logtable0_freq500_uid27
  (input  [7:0] x,
   output [34:0] y);
  wire [34:0] y0;
  wire [34:0] y1;
  wire n2373;
  wire n2376;
  wire n2379;
  wire n2382;
  wire n2385;
  wire n2388;
  wire n2391;
  wire n2394;
  wire n2397;
  wire n2400;
  wire n2403;
  wire n2406;
  wire n2409;
  wire n2412;
  wire n2415;
  wire n2418;
  wire n2421;
  wire n2424;
  wire n2427;
  wire n2430;
  wire n2433;
  wire n2436;
  wire n2439;
  wire n2442;
  wire n2445;
  wire n2448;
  wire n2451;
  wire n2454;
  wire n2457;
  wire n2460;
  wire n2463;
  wire n2466;
  wire n2469;
  wire n2472;
  wire n2475;
  wire n2478;
  wire n2481;
  wire n2484;
  wire n2487;
  wire n2490;
  wire n2493;
  wire n2496;
  wire n2499;
  wire n2502;
  wire n2505;
  wire n2508;
  wire n2511;
  wire n2514;
  wire n2517;
  wire n2520;
  wire n2523;
  wire n2526;
  wire n2529;
  wire n2532;
  wire n2535;
  wire n2538;
  wire n2541;
  wire n2544;
  wire n2547;
  wire n2550;
  wire n2553;
  wire n2556;
  wire n2559;
  wire n2562;
  wire n2565;
  wire n2568;
  wire n2571;
  wire n2574;
  wire n2577;
  wire n2580;
  wire n2583;
  wire n2586;
  wire n2589;
  wire n2592;
  wire n2595;
  wire n2598;
  wire n2601;
  wire n2604;
  wire n2607;
  wire n2610;
  wire n2613;
  wire n2616;
  wire n2619;
  wire n2622;
  wire n2625;
  wire n2628;
  wire n2631;
  wire n2634;
  wire n2637;
  wire n2640;
  wire n2643;
  wire n2646;
  wire n2649;
  wire n2652;
  wire n2655;
  wire n2658;
  wire n2661;
  wire n2664;
  wire n2667;
  wire n2670;
  wire n2673;
  wire n2676;
  wire n2679;
  wire n2682;
  wire n2685;
  wire n2688;
  wire n2691;
  wire n2694;
  wire n2697;
  wire n2700;
  wire n2703;
  wire n2706;
  wire n2709;
  wire n2712;
  wire n2715;
  wire n2718;
  wire n2721;
  wire n2724;
  wire n2727;
  wire n2730;
  wire n2733;
  wire n2736;
  wire n2739;
  wire n2742;
  wire n2745;
  wire n2748;
  wire n2751;
  wire n2754;
  wire n2757;
  wire n2760;
  wire n2763;
  wire n2766;
  wire n2769;
  wire n2772;
  wire n2775;
  wire n2778;
  wire n2781;
  wire n2784;
  wire n2787;
  wire n2790;
  wire n2793;
  wire n2796;
  wire n2799;
  wire n2802;
  wire n2805;
  wire n2808;
  wire n2811;
  wire n2814;
  wire n2817;
  wire n2820;
  wire n2823;
  wire n2826;
  wire n2829;
  wire n2832;
  wire n2835;
  wire n2838;
  wire n2841;
  wire n2844;
  wire n2847;
  wire n2850;
  wire n2853;
  wire n2856;
  wire n2859;
  wire n2862;
  wire n2865;
  wire n2868;
  wire n2871;
  wire n2874;
  wire n2877;
  wire n2880;
  wire n2883;
  wire n2886;
  wire n2889;
  wire n2892;
  wire n2895;
  wire n2898;
  wire n2901;
  wire n2904;
  wire n2907;
  wire n2910;
  wire n2913;
  wire n2916;
  wire n2919;
  wire n2922;
  wire n2925;
  wire n2928;
  wire n2931;
  wire n2934;
  wire n2937;
  wire n2940;
  wire n2943;
  wire n2946;
  wire n2949;
  wire n2952;
  wire n2955;
  wire n2958;
  wire n2961;
  wire n2964;
  wire n2967;
  wire n2970;
  wire n2973;
  wire n2976;
  wire n2979;
  wire n2982;
  wire n2985;
  wire n2988;
  wire n2991;
  wire n2994;
  wire n2997;
  wire n3000;
  wire n3003;
  wire n3006;
  wire n3009;
  wire n3012;
  wire n3015;
  wire n3018;
  wire n3021;
  wire n3024;
  wire n3027;
  wire n3030;
  wire n3033;
  wire n3036;
  wire n3039;
  wire n3042;
  wire n3045;
  wire n3048;
  wire n3051;
  wire n3054;
  wire n3057;
  wire n3060;
  wire n3063;
  wire n3066;
  wire n3069;
  wire n3072;
  wire n3075;
  wire n3078;
  wire n3081;
  wire n3084;
  wire n3087;
  wire n3090;
  wire n3093;
  wire n3096;
  wire n3099;
  wire n3102;
  wire n3105;
  wire n3108;
  wire n3111;
  wire n3114;
  wire n3117;
  wire n3120;
  wire n3123;
  wire n3126;
  wire n3129;
  wire n3132;
  wire n3135;
  wire n3138;
  wire [255:0] n3140;
  reg [34:0] n3141;
  assign y = y1; //(module output)
  /* fppowtf32.vhdl:326:8  */
  assign y0 = n3141; // (signal)
  /* fppowtf32.vhdl:328:8  */
  assign y1 = y0; // (signal)
  /* fppowtf32.vhdl:332:45  */
  assign n2373 = x == 8'b00000000;
  /* fppowtf32.vhdl:333:45  */
  assign n2376 = x == 8'b00000001;
  /* fppowtf32.vhdl:334:45  */
  assign n2379 = x == 8'b00000010;
  /* fppowtf32.vhdl:335:45  */
  assign n2382 = x == 8'b00000011;
  /* fppowtf32.vhdl:336:45  */
  assign n2385 = x == 8'b00000100;
  /* fppowtf32.vhdl:337:45  */
  assign n2388 = x == 8'b00000101;
  /* fppowtf32.vhdl:338:45  */
  assign n2391 = x == 8'b00000110;
  /* fppowtf32.vhdl:339:45  */
  assign n2394 = x == 8'b00000111;
  /* fppowtf32.vhdl:340:45  */
  assign n2397 = x == 8'b00001000;
  /* fppowtf32.vhdl:341:45  */
  assign n2400 = x == 8'b00001001;
  /* fppowtf32.vhdl:342:45  */
  assign n2403 = x == 8'b00001010;
  /* fppowtf32.vhdl:343:45  */
  assign n2406 = x == 8'b00001011;
  /* fppowtf32.vhdl:344:45  */
  assign n2409 = x == 8'b00001100;
  /* fppowtf32.vhdl:345:45  */
  assign n2412 = x == 8'b00001101;
  /* fppowtf32.vhdl:346:45  */
  assign n2415 = x == 8'b00001110;
  /* fppowtf32.vhdl:347:45  */
  assign n2418 = x == 8'b00001111;
  /* fppowtf32.vhdl:348:45  */
  assign n2421 = x == 8'b00010000;
  /* fppowtf32.vhdl:349:45  */
  assign n2424 = x == 8'b00010001;
  /* fppowtf32.vhdl:350:45  */
  assign n2427 = x == 8'b00010010;
  /* fppowtf32.vhdl:351:45  */
  assign n2430 = x == 8'b00010011;
  /* fppowtf32.vhdl:352:45  */
  assign n2433 = x == 8'b00010100;
  /* fppowtf32.vhdl:353:45  */
  assign n2436 = x == 8'b00010101;
  /* fppowtf32.vhdl:354:45  */
  assign n2439 = x == 8'b00010110;
  /* fppowtf32.vhdl:355:45  */
  assign n2442 = x == 8'b00010111;
  /* fppowtf32.vhdl:356:45  */
  assign n2445 = x == 8'b00011000;
  /* fppowtf32.vhdl:357:45  */
  assign n2448 = x == 8'b00011001;
  /* fppowtf32.vhdl:358:45  */
  assign n2451 = x == 8'b00011010;
  /* fppowtf32.vhdl:359:45  */
  assign n2454 = x == 8'b00011011;
  /* fppowtf32.vhdl:360:45  */
  assign n2457 = x == 8'b00011100;
  /* fppowtf32.vhdl:361:45  */
  assign n2460 = x == 8'b00011101;
  /* fppowtf32.vhdl:362:45  */
  assign n2463 = x == 8'b00011110;
  /* fppowtf32.vhdl:363:45  */
  assign n2466 = x == 8'b00011111;
  /* fppowtf32.vhdl:364:45  */
  assign n2469 = x == 8'b00100000;
  /* fppowtf32.vhdl:365:45  */
  assign n2472 = x == 8'b00100001;
  /* fppowtf32.vhdl:366:45  */
  assign n2475 = x == 8'b00100010;
  /* fppowtf32.vhdl:367:45  */
  assign n2478 = x == 8'b00100011;
  /* fppowtf32.vhdl:368:45  */
  assign n2481 = x == 8'b00100100;
  /* fppowtf32.vhdl:369:45  */
  assign n2484 = x == 8'b00100101;
  /* fppowtf32.vhdl:370:45  */
  assign n2487 = x == 8'b00100110;
  /* fppowtf32.vhdl:371:45  */
  assign n2490 = x == 8'b00100111;
  /* fppowtf32.vhdl:372:45  */
  assign n2493 = x == 8'b00101000;
  /* fppowtf32.vhdl:373:45  */
  assign n2496 = x == 8'b00101001;
  /* fppowtf32.vhdl:374:45  */
  assign n2499 = x == 8'b00101010;
  /* fppowtf32.vhdl:375:45  */
  assign n2502 = x == 8'b00101011;
  /* fppowtf32.vhdl:376:45  */
  assign n2505 = x == 8'b00101100;
  /* fppowtf32.vhdl:377:45  */
  assign n2508 = x == 8'b00101101;
  /* fppowtf32.vhdl:378:45  */
  assign n2511 = x == 8'b00101110;
  /* fppowtf32.vhdl:379:45  */
  assign n2514 = x == 8'b00101111;
  /* fppowtf32.vhdl:380:45  */
  assign n2517 = x == 8'b00110000;
  /* fppowtf32.vhdl:381:45  */
  assign n2520 = x == 8'b00110001;
  /* fppowtf32.vhdl:382:45  */
  assign n2523 = x == 8'b00110010;
  /* fppowtf32.vhdl:383:45  */
  assign n2526 = x == 8'b00110011;
  /* fppowtf32.vhdl:384:45  */
  assign n2529 = x == 8'b00110100;
  /* fppowtf32.vhdl:385:45  */
  assign n2532 = x == 8'b00110101;
  /* fppowtf32.vhdl:386:45  */
  assign n2535 = x == 8'b00110110;
  /* fppowtf32.vhdl:387:45  */
  assign n2538 = x == 8'b00110111;
  /* fppowtf32.vhdl:388:45  */
  assign n2541 = x == 8'b00111000;
  /* fppowtf32.vhdl:389:45  */
  assign n2544 = x == 8'b00111001;
  /* fppowtf32.vhdl:390:45  */
  assign n2547 = x == 8'b00111010;
  /* fppowtf32.vhdl:391:45  */
  assign n2550 = x == 8'b00111011;
  /* fppowtf32.vhdl:392:45  */
  assign n2553 = x == 8'b00111100;
  /* fppowtf32.vhdl:393:45  */
  assign n2556 = x == 8'b00111101;
  /* fppowtf32.vhdl:394:45  */
  assign n2559 = x == 8'b00111110;
  /* fppowtf32.vhdl:395:45  */
  assign n2562 = x == 8'b00111111;
  /* fppowtf32.vhdl:396:45  */
  assign n2565 = x == 8'b01000000;
  /* fppowtf32.vhdl:397:45  */
  assign n2568 = x == 8'b01000001;
  /* fppowtf32.vhdl:398:45  */
  assign n2571 = x == 8'b01000010;
  /* fppowtf32.vhdl:399:45  */
  assign n2574 = x == 8'b01000011;
  /* fppowtf32.vhdl:400:45  */
  assign n2577 = x == 8'b01000100;
  /* fppowtf32.vhdl:401:45  */
  assign n2580 = x == 8'b01000101;
  /* fppowtf32.vhdl:402:45  */
  assign n2583 = x == 8'b01000110;
  /* fppowtf32.vhdl:403:45  */
  assign n2586 = x == 8'b01000111;
  /* fppowtf32.vhdl:404:45  */
  assign n2589 = x == 8'b01001000;
  /* fppowtf32.vhdl:405:45  */
  assign n2592 = x == 8'b01001001;
  /* fppowtf32.vhdl:406:45  */
  assign n2595 = x == 8'b01001010;
  /* fppowtf32.vhdl:407:45  */
  assign n2598 = x == 8'b01001011;
  /* fppowtf32.vhdl:408:45  */
  assign n2601 = x == 8'b01001100;
  /* fppowtf32.vhdl:409:45  */
  assign n2604 = x == 8'b01001101;
  /* fppowtf32.vhdl:410:45  */
  assign n2607 = x == 8'b01001110;
  /* fppowtf32.vhdl:411:45  */
  assign n2610 = x == 8'b01001111;
  /* fppowtf32.vhdl:412:45  */
  assign n2613 = x == 8'b01010000;
  /* fppowtf32.vhdl:413:45  */
  assign n2616 = x == 8'b01010001;
  /* fppowtf32.vhdl:414:45  */
  assign n2619 = x == 8'b01010010;
  /* fppowtf32.vhdl:415:45  */
  assign n2622 = x == 8'b01010011;
  /* fppowtf32.vhdl:416:45  */
  assign n2625 = x == 8'b01010100;
  /* fppowtf32.vhdl:417:45  */
  assign n2628 = x == 8'b01010101;
  /* fppowtf32.vhdl:418:45  */
  assign n2631 = x == 8'b01010110;
  /* fppowtf32.vhdl:419:45  */
  assign n2634 = x == 8'b01010111;
  /* fppowtf32.vhdl:420:45  */
  assign n2637 = x == 8'b01011000;
  /* fppowtf32.vhdl:421:45  */
  assign n2640 = x == 8'b01011001;
  /* fppowtf32.vhdl:422:45  */
  assign n2643 = x == 8'b01011010;
  /* fppowtf32.vhdl:423:45  */
  assign n2646 = x == 8'b01011011;
  /* fppowtf32.vhdl:424:45  */
  assign n2649 = x == 8'b01011100;
  /* fppowtf32.vhdl:425:45  */
  assign n2652 = x == 8'b01011101;
  /* fppowtf32.vhdl:426:45  */
  assign n2655 = x == 8'b01011110;
  /* fppowtf32.vhdl:427:45  */
  assign n2658 = x == 8'b01011111;
  /* fppowtf32.vhdl:428:45  */
  assign n2661 = x == 8'b01100000;
  /* fppowtf32.vhdl:429:45  */
  assign n2664 = x == 8'b01100001;
  /* fppowtf32.vhdl:430:45  */
  assign n2667 = x == 8'b01100010;
  /* fppowtf32.vhdl:431:45  */
  assign n2670 = x == 8'b01100011;
  /* fppowtf32.vhdl:432:45  */
  assign n2673 = x == 8'b01100100;
  /* fppowtf32.vhdl:433:45  */
  assign n2676 = x == 8'b01100101;
  /* fppowtf32.vhdl:434:45  */
  assign n2679 = x == 8'b01100110;
  /* fppowtf32.vhdl:435:45  */
  assign n2682 = x == 8'b01100111;
  /* fppowtf32.vhdl:436:45  */
  assign n2685 = x == 8'b01101000;
  /* fppowtf32.vhdl:437:45  */
  assign n2688 = x == 8'b01101001;
  /* fppowtf32.vhdl:438:45  */
  assign n2691 = x == 8'b01101010;
  /* fppowtf32.vhdl:439:45  */
  assign n2694 = x == 8'b01101011;
  /* fppowtf32.vhdl:440:45  */
  assign n2697 = x == 8'b01101100;
  /* fppowtf32.vhdl:441:45  */
  assign n2700 = x == 8'b01101101;
  /* fppowtf32.vhdl:442:45  */
  assign n2703 = x == 8'b01101110;
  /* fppowtf32.vhdl:443:45  */
  assign n2706 = x == 8'b01101111;
  /* fppowtf32.vhdl:444:45  */
  assign n2709 = x == 8'b01110000;
  /* fppowtf32.vhdl:445:45  */
  assign n2712 = x == 8'b01110001;
  /* fppowtf32.vhdl:446:45  */
  assign n2715 = x == 8'b01110010;
  /* fppowtf32.vhdl:447:45  */
  assign n2718 = x == 8'b01110011;
  /* fppowtf32.vhdl:448:45  */
  assign n2721 = x == 8'b01110100;
  /* fppowtf32.vhdl:449:45  */
  assign n2724 = x == 8'b01110101;
  /* fppowtf32.vhdl:450:45  */
  assign n2727 = x == 8'b01110110;
  /* fppowtf32.vhdl:451:45  */
  assign n2730 = x == 8'b01110111;
  /* fppowtf32.vhdl:452:45  */
  assign n2733 = x == 8'b01111000;
  /* fppowtf32.vhdl:453:45  */
  assign n2736 = x == 8'b01111001;
  /* fppowtf32.vhdl:454:45  */
  assign n2739 = x == 8'b01111010;
  /* fppowtf32.vhdl:455:45  */
  assign n2742 = x == 8'b01111011;
  /* fppowtf32.vhdl:456:45  */
  assign n2745 = x == 8'b01111100;
  /* fppowtf32.vhdl:457:45  */
  assign n2748 = x == 8'b01111101;
  /* fppowtf32.vhdl:458:45  */
  assign n2751 = x == 8'b01111110;
  /* fppowtf32.vhdl:459:45  */
  assign n2754 = x == 8'b01111111;
  /* fppowtf32.vhdl:460:45  */
  assign n2757 = x == 8'b10000000;
  /* fppowtf32.vhdl:461:45  */
  assign n2760 = x == 8'b10000001;
  /* fppowtf32.vhdl:462:45  */
  assign n2763 = x == 8'b10000010;
  /* fppowtf32.vhdl:463:45  */
  assign n2766 = x == 8'b10000011;
  /* fppowtf32.vhdl:464:45  */
  assign n2769 = x == 8'b10000100;
  /* fppowtf32.vhdl:465:45  */
  assign n2772 = x == 8'b10000101;
  /* fppowtf32.vhdl:466:45  */
  assign n2775 = x == 8'b10000110;
  /* fppowtf32.vhdl:467:45  */
  assign n2778 = x == 8'b10000111;
  /* fppowtf32.vhdl:468:45  */
  assign n2781 = x == 8'b10001000;
  /* fppowtf32.vhdl:469:45  */
  assign n2784 = x == 8'b10001001;
  /* fppowtf32.vhdl:470:45  */
  assign n2787 = x == 8'b10001010;
  /* fppowtf32.vhdl:471:45  */
  assign n2790 = x == 8'b10001011;
  /* fppowtf32.vhdl:472:45  */
  assign n2793 = x == 8'b10001100;
  /* fppowtf32.vhdl:473:45  */
  assign n2796 = x == 8'b10001101;
  /* fppowtf32.vhdl:474:45  */
  assign n2799 = x == 8'b10001110;
  /* fppowtf32.vhdl:475:45  */
  assign n2802 = x == 8'b10001111;
  /* fppowtf32.vhdl:476:45  */
  assign n2805 = x == 8'b10010000;
  /* fppowtf32.vhdl:477:45  */
  assign n2808 = x == 8'b10010001;
  /* fppowtf32.vhdl:478:45  */
  assign n2811 = x == 8'b10010010;
  /* fppowtf32.vhdl:479:45  */
  assign n2814 = x == 8'b10010011;
  /* fppowtf32.vhdl:480:45  */
  assign n2817 = x == 8'b10010100;
  /* fppowtf32.vhdl:481:45  */
  assign n2820 = x == 8'b10010101;
  /* fppowtf32.vhdl:482:45  */
  assign n2823 = x == 8'b10010110;
  /* fppowtf32.vhdl:483:45  */
  assign n2826 = x == 8'b10010111;
  /* fppowtf32.vhdl:484:45  */
  assign n2829 = x == 8'b10011000;
  /* fppowtf32.vhdl:485:45  */
  assign n2832 = x == 8'b10011001;
  /* fppowtf32.vhdl:486:45  */
  assign n2835 = x == 8'b10011010;
  /* fppowtf32.vhdl:487:45  */
  assign n2838 = x == 8'b10011011;
  /* fppowtf32.vhdl:488:45  */
  assign n2841 = x == 8'b10011100;
  /* fppowtf32.vhdl:489:45  */
  assign n2844 = x == 8'b10011101;
  /* fppowtf32.vhdl:490:45  */
  assign n2847 = x == 8'b10011110;
  /* fppowtf32.vhdl:491:45  */
  assign n2850 = x == 8'b10011111;
  /* fppowtf32.vhdl:492:45  */
  assign n2853 = x == 8'b10100000;
  /* fppowtf32.vhdl:493:45  */
  assign n2856 = x == 8'b10100001;
  /* fppowtf32.vhdl:494:45  */
  assign n2859 = x == 8'b10100010;
  /* fppowtf32.vhdl:495:45  */
  assign n2862 = x == 8'b10100011;
  /* fppowtf32.vhdl:496:45  */
  assign n2865 = x == 8'b10100100;
  /* fppowtf32.vhdl:497:45  */
  assign n2868 = x == 8'b10100101;
  /* fppowtf32.vhdl:498:45  */
  assign n2871 = x == 8'b10100110;
  /* fppowtf32.vhdl:499:45  */
  assign n2874 = x == 8'b10100111;
  /* fppowtf32.vhdl:500:45  */
  assign n2877 = x == 8'b10101000;
  /* fppowtf32.vhdl:501:45  */
  assign n2880 = x == 8'b10101001;
  /* fppowtf32.vhdl:502:45  */
  assign n2883 = x == 8'b10101010;
  /* fppowtf32.vhdl:503:45  */
  assign n2886 = x == 8'b10101011;
  /* fppowtf32.vhdl:504:45  */
  assign n2889 = x == 8'b10101100;
  /* fppowtf32.vhdl:505:45  */
  assign n2892 = x == 8'b10101101;
  /* fppowtf32.vhdl:506:45  */
  assign n2895 = x == 8'b10101110;
  /* fppowtf32.vhdl:507:45  */
  assign n2898 = x == 8'b10101111;
  /* fppowtf32.vhdl:508:45  */
  assign n2901 = x == 8'b10110000;
  /* fppowtf32.vhdl:509:45  */
  assign n2904 = x == 8'b10110001;
  /* fppowtf32.vhdl:510:45  */
  assign n2907 = x == 8'b10110010;
  /* fppowtf32.vhdl:511:45  */
  assign n2910 = x == 8'b10110011;
  /* fppowtf32.vhdl:512:45  */
  assign n2913 = x == 8'b10110100;
  /* fppowtf32.vhdl:513:45  */
  assign n2916 = x == 8'b10110101;
  /* fppowtf32.vhdl:514:45  */
  assign n2919 = x == 8'b10110110;
  /* fppowtf32.vhdl:515:45  */
  assign n2922 = x == 8'b10110111;
  /* fppowtf32.vhdl:516:45  */
  assign n2925 = x == 8'b10111000;
  /* fppowtf32.vhdl:517:45  */
  assign n2928 = x == 8'b10111001;
  /* fppowtf32.vhdl:518:45  */
  assign n2931 = x == 8'b10111010;
  /* fppowtf32.vhdl:519:45  */
  assign n2934 = x == 8'b10111011;
  /* fppowtf32.vhdl:520:45  */
  assign n2937 = x == 8'b10111100;
  /* fppowtf32.vhdl:521:45  */
  assign n2940 = x == 8'b10111101;
  /* fppowtf32.vhdl:522:45  */
  assign n2943 = x == 8'b10111110;
  /* fppowtf32.vhdl:523:45  */
  assign n2946 = x == 8'b10111111;
  /* fppowtf32.vhdl:524:45  */
  assign n2949 = x == 8'b11000000;
  /* fppowtf32.vhdl:525:45  */
  assign n2952 = x == 8'b11000001;
  /* fppowtf32.vhdl:526:45  */
  assign n2955 = x == 8'b11000010;
  /* fppowtf32.vhdl:527:45  */
  assign n2958 = x == 8'b11000011;
  /* fppowtf32.vhdl:528:45  */
  assign n2961 = x == 8'b11000100;
  /* fppowtf32.vhdl:529:45  */
  assign n2964 = x == 8'b11000101;
  /* fppowtf32.vhdl:530:45  */
  assign n2967 = x == 8'b11000110;
  /* fppowtf32.vhdl:531:45  */
  assign n2970 = x == 8'b11000111;
  /* fppowtf32.vhdl:532:45  */
  assign n2973 = x == 8'b11001000;
  /* fppowtf32.vhdl:533:45  */
  assign n2976 = x == 8'b11001001;
  /* fppowtf32.vhdl:534:45  */
  assign n2979 = x == 8'b11001010;
  /* fppowtf32.vhdl:535:45  */
  assign n2982 = x == 8'b11001011;
  /* fppowtf32.vhdl:536:45  */
  assign n2985 = x == 8'b11001100;
  /* fppowtf32.vhdl:537:45  */
  assign n2988 = x == 8'b11001101;
  /* fppowtf32.vhdl:538:45  */
  assign n2991 = x == 8'b11001110;
  /* fppowtf32.vhdl:539:45  */
  assign n2994 = x == 8'b11001111;
  /* fppowtf32.vhdl:540:45  */
  assign n2997 = x == 8'b11010000;
  /* fppowtf32.vhdl:541:45  */
  assign n3000 = x == 8'b11010001;
  /* fppowtf32.vhdl:542:45  */
  assign n3003 = x == 8'b11010010;
  /* fppowtf32.vhdl:543:45  */
  assign n3006 = x == 8'b11010011;
  /* fppowtf32.vhdl:544:45  */
  assign n3009 = x == 8'b11010100;
  /* fppowtf32.vhdl:545:45  */
  assign n3012 = x == 8'b11010101;
  /* fppowtf32.vhdl:546:45  */
  assign n3015 = x == 8'b11010110;
  /* fppowtf32.vhdl:547:45  */
  assign n3018 = x == 8'b11010111;
  /* fppowtf32.vhdl:548:45  */
  assign n3021 = x == 8'b11011000;
  /* fppowtf32.vhdl:549:45  */
  assign n3024 = x == 8'b11011001;
  /* fppowtf32.vhdl:550:45  */
  assign n3027 = x == 8'b11011010;
  /* fppowtf32.vhdl:551:45  */
  assign n3030 = x == 8'b11011011;
  /* fppowtf32.vhdl:552:45  */
  assign n3033 = x == 8'b11011100;
  /* fppowtf32.vhdl:553:45  */
  assign n3036 = x == 8'b11011101;
  /* fppowtf32.vhdl:554:45  */
  assign n3039 = x == 8'b11011110;
  /* fppowtf32.vhdl:555:45  */
  assign n3042 = x == 8'b11011111;
  /* fppowtf32.vhdl:556:45  */
  assign n3045 = x == 8'b11100000;
  /* fppowtf32.vhdl:557:45  */
  assign n3048 = x == 8'b11100001;
  /* fppowtf32.vhdl:558:45  */
  assign n3051 = x == 8'b11100010;
  /* fppowtf32.vhdl:559:45  */
  assign n3054 = x == 8'b11100011;
  /* fppowtf32.vhdl:560:45  */
  assign n3057 = x == 8'b11100100;
  /* fppowtf32.vhdl:561:45  */
  assign n3060 = x == 8'b11100101;
  /* fppowtf32.vhdl:562:45  */
  assign n3063 = x == 8'b11100110;
  /* fppowtf32.vhdl:563:45  */
  assign n3066 = x == 8'b11100111;
  /* fppowtf32.vhdl:564:45  */
  assign n3069 = x == 8'b11101000;
  /* fppowtf32.vhdl:565:45  */
  assign n3072 = x == 8'b11101001;
  /* fppowtf32.vhdl:566:45  */
  assign n3075 = x == 8'b11101010;
  /* fppowtf32.vhdl:567:45  */
  assign n3078 = x == 8'b11101011;
  /* fppowtf32.vhdl:568:45  */
  assign n3081 = x == 8'b11101100;
  /* fppowtf32.vhdl:569:45  */
  assign n3084 = x == 8'b11101101;
  /* fppowtf32.vhdl:570:45  */
  assign n3087 = x == 8'b11101110;
  /* fppowtf32.vhdl:571:45  */
  assign n3090 = x == 8'b11101111;
  /* fppowtf32.vhdl:572:45  */
  assign n3093 = x == 8'b11110000;
  /* fppowtf32.vhdl:573:45  */
  assign n3096 = x == 8'b11110001;
  /* fppowtf32.vhdl:574:45  */
  assign n3099 = x == 8'b11110010;
  /* fppowtf32.vhdl:575:45  */
  assign n3102 = x == 8'b11110011;
  /* fppowtf32.vhdl:576:45  */
  assign n3105 = x == 8'b11110100;
  /* fppowtf32.vhdl:577:45  */
  assign n3108 = x == 8'b11110101;
  /* fppowtf32.vhdl:578:45  */
  assign n3111 = x == 8'b11110110;
  /* fppowtf32.vhdl:579:45  */
  assign n3114 = x == 8'b11110111;
  /* fppowtf32.vhdl:580:45  */
  assign n3117 = x == 8'b11111000;
  /* fppowtf32.vhdl:581:45  */
  assign n3120 = x == 8'b11111001;
  /* fppowtf32.vhdl:582:45  */
  assign n3123 = x == 8'b11111010;
  /* fppowtf32.vhdl:583:45  */
  assign n3126 = x == 8'b11111011;
  /* fppowtf32.vhdl:584:45  */
  assign n3129 = x == 8'b11111100;
  /* fppowtf32.vhdl:585:45  */
  assign n3132 = x == 8'b11111101;
  /* fppowtf32.vhdl:586:45  */
  assign n3135 = x == 8'b11111110;
  /* fppowtf32.vhdl:587:45  */
  assign n3138 = x == 8'b11111111;
  assign n3140 = {n3138, n3135, n3132, n3129, n3126, n3123, n3120, n3117, n3114, n3111, n3108, n3105, n3102, n3099, n3096, n3093, n3090, n3087, n3084, n3081, n3078, n3075, n3072, n3069, n3066, n3063, n3060, n3057, n3054, n3051, n3048, n3045, n3042, n3039, n3036, n3033, n3030, n3027, n3024, n3021, n3018, n3015, n3012, n3009, n3006, n3003, n3000, n2997, n2994, n2991, n2988, n2985, n2982, n2979, n2976, n2973, n2970, n2967, n2964, n2961, n2958, n2955, n2952, n2949, n2946, n2943, n2940, n2937, n2934, n2931, n2928, n2925, n2922, n2919, n2916, n2913, n2910, n2907, n2904, n2901, n2898, n2895, n2892, n2889, n2886, n2883, n2880, n2877, n2874, n2871, n2868, n2865, n2862, n2859, n2856, n2853, n2850, n2847, n2844, n2841, n2838, n2835, n2832, n2829, n2826, n2823, n2820, n2817, n2814, n2811, n2808, n2805, n2802, n2799, n2796, n2793, n2790, n2787, n2784, n2781, n2778, n2775, n2772, n2769, n2766, n2763, n2760, n2757, n2754, n2751, n2748, n2745, n2742, n2739, n2736, n2733, n2730, n2727, n2724, n2721, n2718, n2715, n2712, n2709, n2706, n2703, n2700, n2697, n2694, n2691, n2688, n2685, n2682, n2679, n2676, n2673, n2670, n2667, n2664, n2661, n2658, n2655, n2652, n2649, n2646, n2643, n2640, n2637, n2634, n2631, n2628, n2625, n2622, n2619, n2616, n2613, n2610, n2607, n2604, n2601, n2598, n2595, n2592, n2589, n2586, n2583, n2580, n2577, n2574, n2571, n2568, n2565, n2562, n2559, n2556, n2553, n2550, n2547, n2544, n2541, n2538, n2535, n2532, n2529, n2526, n2523, n2520, n2517, n2514, n2511, n2508, n2505, n2502, n2499, n2496, n2493, n2490, n2487, n2484, n2481, n2478, n2475, n2472, n2469, n2466, n2463, n2460, n2457, n2454, n2451, n2448, n2445, n2442, n2439, n2436, n2433, n2430, n2427, n2424, n2421, n2418, n2415, n2412, n2409, n2406, n2403, n2400, n2397, n2394, n2391, n2388, n2385, n2382, n2379, n2376, n2373};
  /* fppowtf32.vhdl:331:4  */
  always @*
    case (n3140)
      256'b1000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3141 = 35'b11111110111100000111111110101010111;
      256'b0100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3141 = 35'b11111101111100011111110101011001010;
      256'b0010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3141 = 35'b11111101111100011111110101011001010;
      256'b0001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3141 = 35'b11111100111101000111011100010100000;
      256'b0000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3141 = 35'b11111100111101000111011100010100000;
      256'b0000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3141 = 35'b11111011111101111110101011101001111;
      256'b0000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3141 = 35'b11111011111101111110101011101001111;
      256'b0000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3141 = 35'b11111010111111000101011011101111001;
      256'b0000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3141 = 35'b11111010111111000101011011101111001;
      256'b0000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3141 = 35'b11111010000000011011100100111110000;
      256'b0000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3141 = 35'b11111010000000011011100100111110000;
      256'b0000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3141 = 35'b11111001000010000000111111110110001;
      256'b0000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3141 = 35'b11111001000010000000111111110110001;
      256'b0000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3141 = 35'b11111000000011110101100100111100011;
      256'b0000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3141 = 35'b11111000000011110101100100111100011;
      256'b0000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3141 = 35'b11110111000101111001001100111011011;
      256'b0000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3141 = 35'b11110111000101111001001100111011011;
      256'b0000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3141 = 35'b11110110001000001011110000100011000;
      256'b0000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3141 = 35'b11110110001000001011110000100011000;
      256'b0000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3141 = 35'b11110101001010101101001000101000001;
      256'b0000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3141 = 35'b11110101001010101101001000101000001;
      256'b0000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3141 = 35'b11110100001101011101001110000100111;
      256'b0000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3141 = 35'b11110011010000011011111001111000101;
      256'b0000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3141 = 35'b11110011010000011011111001111000101;
      256'b0000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3141 = 35'b11110010010011101001000101000111100;
      256'b0000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3141 = 35'b11110010010011101001000101000111100;
      256'b0000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3141 = 35'b11110001010111000100101000111010101;
      256'b0000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3141 = 35'b11110001010111000100101000111010101;
      256'b0000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3141 = 35'b11110000011010101110011110100000000;
      256'b0000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3141 = 35'b11110000011010101110011110100000000;
      256'b0000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3141 = 35'b11101111011110100110011111001010011;
      256'b0000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3141 = 35'b11101110100010101100100100010001011;
      256'b0000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3141 = 35'b11101110100010101100100100010001011;
      256'b0000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3141 = 35'b11101101100111000000100111010001000;
      256'b0000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3141 = 35'b11101101100111000000100111010001000;
      256'b0000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3141 = 35'b11101100101011100010100001101001111;
      256'b0000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3141 = 35'b11101100101011100010100001101001111;
      256'b0000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3141 = 35'b11101011110000010010001101000001011;
      256'b0000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3141 = 35'b11101010110101001111100011000001000;
      256'b0000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3141 = 35'b11101010110101001111100011000001000;
      256'b0000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3141 = 35'b11101001111010011010011101010110110;
      256'b0000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3141 = 35'b11101001111010011010011101010110110;
      256'b0000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3141 = 35'b11101000111111110010110101110101001;
      256'b0000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3141 = 35'b11101000000101011000100110010010100;
      256'b0000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3141 = 35'b11101000000101011000100110010010100;
      256'b0000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3141 = 35'b11100111001011001011101000101001110;
      256'b0000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3141 = 35'b11100111001011001011101000101001110;
      256'b0000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3141 = 35'b11100110010001001011110110111001111;
      256'b0000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3141 = 35'b11100101010111011001001011000101110;
      256'b0000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3141 = 35'b11100101010111011001001011000101110;
      256'b0000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3141 = 35'b11100100011101110011011111010100010;
      256'b0000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3141 = 35'b11100100011101110011011111010100010;
      256'b0000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3141 = 35'b11100011100100011010101101110000101;
      256'b0000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3141 = 35'b11100010101011001110110000101001101;
      256'b0000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3141 = 35'b11100010101011001110110000101001101;
      256'b0000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3141 = 35'b11100001110010001111100010010001111;
      256'b0000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3141 = 35'b11100000111001011100111101000000000;
      256'b0000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3141 = 35'b11100000111001011100111101000000000;
      256'b0000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3141 = 35'b11100000000000110110111011001110001;
      256'b0000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3141 = 35'b11100000000000110110111011001110001;
      256'b0000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3141 = 35'b11011111001000011101010111011010011;
      256'b0000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3141 = 35'b11011110010000010000001100000110011;
      256'b0000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3141 = 35'b11011110010000010000001100000110011;
      256'b0000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3141 = 35'b11011101011000001111010011110111010;
      256'b0000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3141 = 35'b11011100100000011010101001010101101;
      256'b0000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3141 = 35'b11011100100000011010101001010101101;
      256'b0000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3141 = 35'b11011011101000110010000111001101111;
      256'b0000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3141 = 35'b11011010110001010101101000001111110;
      256'b0000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3141 = 35'b11011010110001010101101000001111110;
      256'b0000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3141 = 35'b11011001111010000101000111001110010;
      256'b0000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3141 = 35'b11011001000011000000011110111111110;
      256'b0000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3141 = 35'b11011001000011000000011110111111110;
      256'b0000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3141 = 35'b11011000001100000111101010011110001;
      256'b0000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3141 = 35'b11010111010101011010100100100110011;
      256'b0000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3141 = 35'b11010111010101011010100100100110011;
      256'b0000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3141 = 35'b11010110011110111001001000011000110;
      256'b0000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3141 = 35'b11010101101000100011010000111000110;
      256'b0000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3141 = 35'b11010100110010011000111001001100110;
      256'b0000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3141 = 35'b11010100110010011000111001001100110;
      256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3141 = 35'b11010011111100011001111100011110110;
      256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3141 = 35'b11010011000110100110010101111011001;
      256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3141 = 35'b11010011000110100110010101111011001;
      256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3141 = 35'b11010010010000111110000000110001110;
      256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3141 = 35'b11010001011011100000111000010101100;
      256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3141 = 35'b11010001011011100000111000010101100;
      256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3141 = 35'b11010000100110001110110111111011111;
      256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3141 = 35'b11001111110001000111111010111101100;
      256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3141 = 35'b11001110111100001011111100110101110;
      256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3141 = 35'b11001110111100001011111100110101110;
      256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3141 = 35'b11001110000111011010111001000011000;
      256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3141 = 35'b11001101010010110100101011000110001;
      256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3141 = 35'b11001100011110011001001110100011000;
      256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3141 = 35'b11001100011110011001001110100011000;
      256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3141 = 35'b11001011101010001000011111000000010;
      256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3141 = 35'b11001010110110000010011000000111000;
      256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3141 = 35'b11001010000010000110110101100011000;
      256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3141 = 35'b11001010000010000110110101100011000;
      256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3141 = 35'b11001001001110010101110011000010111;
      256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3141 = 35'b11001000011010101111001100010111101;
      256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3141 = 35'b11000111100111010010111101010100111;
      256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3141 = 35'b11000111100111010010111101010100111;
      256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3141 = 35'b11000110110100000001000001110000110;
      256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3141 = 35'b11000110000000111001010101100100000;
      256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3141 = 35'b11000101001101111011110100101001011;
      256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3141 = 35'b11000100011011001000011010111110101;
      256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3141 = 35'b11000100011011001000011010111110101;
      256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3141 = 35'b11000011101000011111000100100011101;
      256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3141 = 35'b11000010110101111111101101011010101;
      256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3141 = 35'b11000010000011101010010001101000010;
      256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3141 = 35'b11000001010001011110101101010011011;
      256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3141 = 35'b11000001010001011110101101010011011;
      256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3141 = 35'b11000000011111011100111100100101010;
      256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3141 = 35'b10111111101101100100111011101001010;
      256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3141 = 35'b10111110111011110110100110101101010;
      256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3141 = 35'b10111110001010010001111010000000110;
      256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3141 = 35'b10111110001010010001111010000000110;
      256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3141 = 35'b10111101011000110110110001110110010;
      256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3141 = 35'b10111100100111100101001010100001100;
      256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3141 = 35'b10111011110110011101000000011001010;
      256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3141 = 35'b10111011000101011110001111110101110;
      256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3141 = 35'b10111010010100101000110101010001010;
      256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3141 = 35'b10111001100011111100101101001000110;
      256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3141 = 35'b10111001100011111100101101001000110;
      256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3141 = 35'b10111000110011011001110011111010011;
      256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3141 = 35'b10111000000011000000000110000110111;
      256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3141 = 35'b10110111010010101111100000010000110;
      256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3141 = 35'b10110110100010100111111110111100100;
      256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3141 = 35'b10110101110010101001011110110000100;
      256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3141 = 35'b01100101101111101000110100001100010;
      256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3141 = 35'b01100101101111101000110100001100010;
      256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3141 = 35'b01100100010000101010000110001101100;
      256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3141 = 35'b01100100010000101010000110001101100;
      256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3141 = 35'b01100100010000101010000110001101100;
      256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3141 = 35'b01100010110010001110011010100010010;
      256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3141 = 35'b01100010110010001110011010100010010;
      256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3141 = 35'b01100001010100010101010111011101110;
      256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3141 = 35'b01100001010100010101010111011101110;
      256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3141 = 35'b01011111110110111110100011101111011;
      256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3141 = 35'b01011111110110111110100011101111011;
      256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3141 = 35'b01011110011010001001100110100010000;
      256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3141 = 35'b01011110011010001001100110100010000;
      256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3141 = 35'b01011100111101110110000111011011001;
      256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3141 = 35'b01011100111101110110000111011011001;
      256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3141 = 35'b01011011100010000011101110011010110;
      256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3141 = 35'b01011011100010000011101110011010110;
      256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3141 = 35'b01011010000110110010000011111010100;
      256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3141 = 35'b01011010000110110010000011111010100;
      256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3141 = 35'b01011000101100000000110000101101000;
      256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3141 = 35'b01011000101100000000110000101101000;
      256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3141 = 35'b01010111010001101111011101111101011;
      256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3141 = 35'b01010111010001101111011101111101011;
      256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3141 = 35'b01010101110111111101110101001111001;
      256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3141 = 35'b01010101110111111101110101001111001;
      256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3141 = 35'b01010100011110101011100000011100111;
      256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3141 = 35'b01010100011110101011100000011100111;
      256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3141 = 35'b01010011000101111000001001111000011;
      256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3141 = 35'b01010011000101111000001001111000011;
      256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3141 = 35'b01010001101101100011011100001001110;
      256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3141 = 35'b01010001101101100011011100001001110;
      256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3141 = 35'b01010000010101101101000010001111010;
      256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3141 = 35'b01010000010101101101000010001111010;
      256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3141 = 35'b01001110111110010100100111011100110;
      256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3141 = 35'b01001110111110010100100111011100110;
      256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3141 = 35'b01001101100111011001110111011011000;
      256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3141 = 35'b01001101100111011001110111011011000;
      256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3141 = 35'b01001100010000111100011110000111010;
      256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3141 = 35'b01001100010000111100011110000111010;
      256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3141 = 35'b01001010111010111100000111110011100;
      256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3141 = 35'b01001001100101011000100001000100110;
      256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3141 = 35'b01001001100101011000100001000100110;
      256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3141 = 35'b01001000010000010001010110110100010;
      256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3141 = 35'b01001000010000010001010110110100010;
      256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3141 = 35'b01000110111011100110010110001101100;
      256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3141 = 35'b01000110111011100110010110001101100;
      256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000: n3141 = 35'b01000101100111010111001100101110110;
      256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000: n3141 = 35'b01000100010011100011101000001000101;
      256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000: n3141 = 35'b01000100010011100011101000001000101;
      256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000: n3141 = 35'b01000011000000001011010110011101100;
      256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000: n3141 = 35'b01000011000000001011010110011101100;
      256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000: n3141 = 35'b01000001101101001110000110000001010;
      256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000: n3141 = 35'b01000001101101001110000110000001010;
      256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000: n3141 = 35'b01000000011010101011100101011000101;
      256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000: n3141 = 35'b00111111001000100011100011011001011;
      256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000: n3141 = 35'b00111111001000100011100011011001011;
      256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000: n3141 = 35'b00111101110110110101101111001001110;
      256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000: n3141 = 35'b00111100100101100001110111111111110;
      256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000: n3141 = 35'b00111100100101100001110111111111110;
      256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000: n3141 = 35'b00111011010100100111101101100001101;
      256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000: n3141 = 35'b00111011010100100111101101100001101;
      256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000: n3141 = 35'b00111010000100000110111111100100110;
      256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000: n3141 = 35'b00111000110011111111011110001101111;
      256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000: n3141 = 35'b00111000110011111111011110001101111;
      256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000: n3141 = 35'b00110111100100010000111001110000100;
      256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000: n3141 = 35'b00110110010100111011000010101110110;
      256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000: n3141 = 35'b00110110010100111011000010101110110;
      256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000: n3141 = 35'b00110101000101111101101001111001001;
      256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000: n3141 = 35'b00110011110111011000100000001110000;
      256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000: n3141 = 35'b00110011110111011000100000001110000;
      256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000: n3141 = 35'b00110010101001001011010110111010000;
      256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000: n3141 = 35'b00110001011011010101111111010110100;
      256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000: n3141 = 35'b00110001011011010101111111010110100;
      256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000: n3141 = 35'b00110000001101111000001011001010101;
      256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000: n3141 = 35'b00101111000000110001101100001010100;
      256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000: n3141 = 35'b00101111000000110001101100001010100;
      256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000: n3141 = 35'b00101101110100000010010100010110111;
      256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000: n3141 = 35'b00101100100111101001110101111101001;
      256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000: n3141 = 35'b00101100100111101001110101111101001;
      256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000: n3141 = 35'b00101011011011101000000011010110101;
      256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000: n3141 = 35'b00101010001111111100101111001001010;
      256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000: n3141 = 35'b00101001000100100111101100000110011;
      256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000: n3141 = 35'b00101001000100100111101100000110011;
      256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000: n3141 = 35'b00100111111001101000101101001011010;
      256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000: n3141 = 35'b00100110101110111111100101100000001;
      256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000: n3141 = 35'b00100110101110111111100101100000001;
      256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000: n3141 = 35'b00100101100100101100001000011001000;
      256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000: n3141 = 35'b00100100011010101110001001010100100;
      256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000: n3141 = 35'b00100011010001000101011011111100010;
      256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000: n3141 = 35'b00100011010001000101011011111100010;
      256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000: n3141 = 35'b00100010000111110001110100000100010;
      256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000: n3141 = 35'b00100000111110110011000101101011010;
      256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000: n3141 = 35'b00011111110110001001000100111001111;
      256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000: n3141 = 35'b00011111110110001001000100111001111;
      256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000: n3141 = 35'b00011110101101110011100110000011000;
      256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000: n3141 = 35'b00011101100101110010011101100011100;
      256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000: n3141 = 35'b00011100011110000101100000000001110;
      256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000: n3141 = 35'b00011011010110101100100010001101101;
      256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000: n3141 = 35'b00011011010110101100100010001101101;
      256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000: n3141 = 35'b00011010001111100111011001000000110;
      256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000: n3141 = 35'b00011001001000110101111001011101011;
      256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000: n3141 = 35'b00011000000010010111111000101111010;
      256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000: n3141 = 35'b00010110111100001101001100001010111;
      256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000: n3141 = 35'b00010101110110010101101001001101101;
      256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000: n3141 = 35'b00010101110110010101101001001101101;
      256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000: n3141 = 35'b00010100110000110001000101011101001;
      256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000: n3141 = 35'b00010011101011011111010110100111110;
      256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000: n3141 = 35'b00010010100110100000010010100100010;
      256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000: n3141 = 35'b00010001100001110011101111010001010;
      256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000: n3141 = 35'b00010000011101011001100010110101101;
      256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000: n3141 = 35'b00001111011001010001100011100000000;
      256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000: n3141 = 35'b00001111011001010001100011100000000;
      256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000: n3141 = 35'b00001110010101011011100111100110111;
      256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000: n3141 = 35'b00001101010001110111100101101000100;
      256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000: n3141 = 35'b00001100001110100101010100001010010;
      256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000: n3141 = 35'b00001011001011100100101001111001011;
      256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000: n3141 = 35'b00001010001000110101011101101010001;
      256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000: n3141 = 35'b00001001000110010111100110010111110;
      256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000: n3141 = 35'b00001000000100001010111011000101000;
      256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000: n3141 = 35'b00000111000010001111010010111011000;
      256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000: n3141 = 35'b00000110000000100100100101001010010;
      256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000: n3141 = 35'b00000100111111001010101001001001011;
      256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000: n3141 = 35'b00000011111110000001010110010110001;
      256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000: n3141 = 35'b00000010111101001000100100010100100;
      256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000: n3141 = 35'b00000001111100100000001010101110110;
      256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100: n3141 = 35'b00000000111100001000000001010101101;
      256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010: n3141 = 35'b11111111111100000000000000000000000;
      256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001: n3141 = 35'b11111111111100000000000000000000000;
      default: n3141 = 35'bX;
    endcase
endmodule

module intadder_24_freq500_uid25
  (input  clk,
   input  [23:0] x,
   input  [23:0] y,
   input  cin,
   output [23:0] r);
  wire [23:0] rtmp;
  wire [23:0] x_d1;
  wire [23:0] x_d2;
  wire [23:0] x_d3;
  wire [23:0] y_d1;
  wire cin_d1;
  wire cin_d2;
  wire cin_d3;
  wire cin_d4;
  wire cin_d5;
  wire cin_d6;
  wire [23:0] n2357;
  wire [23:0] n2358;
  wire [23:0] n2359;
  reg [23:0] n2360;
  reg [23:0] n2361;
  reg [23:0] n2362;
  reg [23:0] n2363;
  reg n2364;
  reg n2365;
  reg n2366;
  reg n2367;
  reg n2368;
  reg n2369;
  assign r = rtmp; //(module output)
  /* fppowtf32.vhdl:2618:8  */
  assign rtmp = n2359; // (signal)
  /* fppowtf32.vhdl:2620:8  */
  assign x_d1 = n2360; // (signal)
  /* fppowtf32.vhdl:2620:14  */
  assign x_d2 = n2361; // (signal)
  /* fppowtf32.vhdl:2620:20  */
  assign x_d3 = n2362; // (signal)
  /* fppowtf32.vhdl:2622:8  */
  assign y_d1 = n2363; // (signal)
  /* fppowtf32.vhdl:2624:8  */
  assign cin_d1 = n2364; // (signal)
  /* fppowtf32.vhdl:2624:16  */
  assign cin_d2 = n2365; // (signal)
  /* fppowtf32.vhdl:2624:24  */
  assign cin_d3 = n2366; // (signal)
  /* fppowtf32.vhdl:2624:32  */
  assign cin_d4 = n2367; // (signal)
  /* fppowtf32.vhdl:2624:40  */
  assign cin_d5 = n2368; // (signal)
  /* fppowtf32.vhdl:2624:48  */
  assign cin_d6 = n2369; // (signal)
  /* fppowtf32.vhdl:2642:17  */
  assign n2357 = x_d3 + y_d1;
  /* fppowtf32.vhdl:2642:24  */
  assign n2358 = {23'b0, cin_d6};  //  uext
  /* fppowtf32.vhdl:2642:24  */
  assign n2359 = n2357 + n2358;
  /* fppowtf32.vhdl:2629:10  */
  always @(posedge clk)
    n2360 <= x;
  /* fppowtf32.vhdl:2629:10  */
  always @(posedge clk)
    n2361 <= x_d1;
  /* fppowtf32.vhdl:2629:10  */
  always @(posedge clk)
    n2362 <= x_d2;
  /* fppowtf32.vhdl:2629:10  */
  always @(posedge clk)
    n2363 <= y;
  /* fppowtf32.vhdl:2629:10  */
  always @(posedge clk)
    n2364 <= cin;
  /* fppowtf32.vhdl:2629:10  */
  always @(posedge clk)
    n2365 <= cin_d1;
  /* fppowtf32.vhdl:2629:10  */
  always @(posedge clk)
    n2366 <= cin_d2;
  /* fppowtf32.vhdl:2629:10  */
  always @(posedge clk)
    n2367 <= cin_d3;
  /* fppowtf32.vhdl:2629:10  */
  always @(posedge clk)
    n2368 <= cin_d4;
  /* fppowtf32.vhdl:2629:10  */
  always @(posedge clk)
    n2369 <= cin_d5;
endmodule

module intadder_24_freq500_uid22
  (input  clk,
   input  [23:0] x,
   input  [23:0] y,
   input  cin,
   output [23:0] r);
  wire cin_1;
  wire cin_1_d1;
  wire cin_1_d2;
  wire cin_1_d3;
  wire [24:0] x_1;
  wire [24:0] x_1_d1;
  wire [24:0] y_1;
  wire [24:0] y_1_d1;
  wire [24:0] s_1;
  wire [23:0] r_1;
  wire [24:0] n2330;
  wire [24:0] n2332;
  wire [24:0] n2333;
  wire [24:0] n2334;
  wire [24:0] n2335;
  wire [23:0] n2336;
  reg n2337;
  reg n2338;
  reg n2339;
  reg [24:0] n2340;
  reg [24:0] n2341;
  assign r = r_1; //(module output)
  /* fppowtf32.vhdl:2557:15  */
  assign cin_1_d1 = n2337; // (signal)
  /* fppowtf32.vhdl:2557:25  */
  assign cin_1_d2 = n2338; // (signal)
  /* fppowtf32.vhdl:2557:35  */
  assign cin_1_d3 = n2339; // (signal)
  /* fppowtf32.vhdl:2559:8  */
  assign x_1 = n2330; // (signal)
  /* fppowtf32.vhdl:2559:13  */
  assign x_1_d1 = n2340; // (signal)
  /* fppowtf32.vhdl:2561:8  */
  assign y_1 = n2332; // (signal)
  /* fppowtf32.vhdl:2561:13  */
  assign y_1_d1 = n2341; // (signal)
  /* fppowtf32.vhdl:2563:8  */
  assign s_1 = n2335; // (signal)
  /* fppowtf32.vhdl:2565:8  */
  assign r_1 = n2336; // (signal)
  /* fppowtf32.vhdl:2579:15  */
  assign n2330 = {1'b0, x};
  /* fppowtf32.vhdl:2580:15  */
  assign n2332 = {1'b0, y};
  /* fppowtf32.vhdl:2581:18  */
  assign n2333 = x_1_d1 + y_1_d1;
  /* fppowtf32.vhdl:2581:27  */
  assign n2334 = {24'b0, cin_1_d3};  //  uext
  /* fppowtf32.vhdl:2581:27  */
  assign n2335 = n2333 + n2334;
  /* fppowtf32.vhdl:2582:14  */
  assign n2336 = s_1[23:0]; // extract
  /* fppowtf32.vhdl:2570:10  */
  always @(posedge clk)
    n2337 <= cin_1;
  /* fppowtf32.vhdl:2570:10  */
  always @(posedge clk)
    n2338 <= cin_1_d1;
  /* fppowtf32.vhdl:2570:10  */
  always @(posedge clk)
    n2339 <= cin_1_d2;
  /* fppowtf32.vhdl:2570:10  */
  always @(posedge clk)
    n2340 <= x_1;
  /* fppowtf32.vhdl:2570:10  */
  always @(posedge clk)
    n2341 <= y_1;
endmodule

module intadder_24_freq500_uid19
  (input  clk,
   input  [23:0] x,
   input  [23:0] y,
   input  cin,
   output [23:0] r);
  wire cin_1;
  wire cin_1_d1;
  wire cin_1_d2;
  wire [24:0] x_1;
  wire [24:0] x_1_d1;
  wire [24:0] y_1;
  wire [24:0] y_1_d1;
  wire [24:0] s_1;
  wire [23:0] r_1;
  wire [24:0] n2308;
  wire [24:0] n2310;
  wire [24:0] n2311;
  wire [24:0] n2312;
  wire [24:0] n2313;
  wire [23:0] n2314;
  reg n2315;
  reg n2316;
  reg [24:0] n2317;
  reg [24:0] n2318;
  assign r = r_1; //(module output)
  /* fppowtf32.vhdl:2497:15  */
  assign cin_1_d1 = n2315; // (signal)
  /* fppowtf32.vhdl:2497:25  */
  assign cin_1_d2 = n2316; // (signal)
  /* fppowtf32.vhdl:2499:8  */
  assign x_1 = n2308; // (signal)
  /* fppowtf32.vhdl:2499:13  */
  assign x_1_d1 = n2317; // (signal)
  /* fppowtf32.vhdl:2501:8  */
  assign y_1 = n2310; // (signal)
  /* fppowtf32.vhdl:2501:13  */
  assign y_1_d1 = n2318; // (signal)
  /* fppowtf32.vhdl:2503:8  */
  assign s_1 = n2313; // (signal)
  /* fppowtf32.vhdl:2505:8  */
  assign r_1 = n2314; // (signal)
  /* fppowtf32.vhdl:2518:15  */
  assign n2308 = {1'b0, x};
  /* fppowtf32.vhdl:2519:15  */
  assign n2310 = {1'b0, y};
  /* fppowtf32.vhdl:2520:18  */
  assign n2311 = x_1_d1 + y_1_d1;
  /* fppowtf32.vhdl:2520:27  */
  assign n2312 = {24'b0, cin_1_d2};  //  uext
  /* fppowtf32.vhdl:2520:27  */
  assign n2313 = n2311 + n2312;
  /* fppowtf32.vhdl:2521:14  */
  assign n2314 = s_1[23:0]; // extract
  /* fppowtf32.vhdl:2510:10  */
  always @(posedge clk)
    n2315 <= cin_1;
  /* fppowtf32.vhdl:2510:10  */
  always @(posedge clk)
    n2316 <= cin_1_d1;
  /* fppowtf32.vhdl:2510:10  */
  always @(posedge clk)
    n2317 <= x_1;
  /* fppowtf32.vhdl:2510:10  */
  always @(posedge clk)
    n2318 <= y_1;
endmodule

module inva0table_freq500_uid15
  (input  [7:0] x,
   output [8:0] y);
  wire [8:0] y0;
  wire [8:0] y1;
  wire n1529;
  wire n1532;
  wire n1535;
  wire n1538;
  wire n1541;
  wire n1544;
  wire n1547;
  wire n1550;
  wire n1553;
  wire n1556;
  wire n1559;
  wire n1562;
  wire n1565;
  wire n1568;
  wire n1571;
  wire n1574;
  wire n1577;
  wire n1580;
  wire n1583;
  wire n1586;
  wire n1589;
  wire n1592;
  wire n1595;
  wire n1598;
  wire n1601;
  wire n1604;
  wire n1607;
  wire n1610;
  wire n1613;
  wire n1616;
  wire n1619;
  wire n1622;
  wire n1625;
  wire n1628;
  wire n1631;
  wire n1634;
  wire n1637;
  wire n1640;
  wire n1643;
  wire n1646;
  wire n1649;
  wire n1652;
  wire n1655;
  wire n1658;
  wire n1661;
  wire n1664;
  wire n1667;
  wire n1670;
  wire n1673;
  wire n1676;
  wire n1679;
  wire n1682;
  wire n1685;
  wire n1688;
  wire n1691;
  wire n1694;
  wire n1697;
  wire n1700;
  wire n1703;
  wire n1706;
  wire n1709;
  wire n1712;
  wire n1715;
  wire n1718;
  wire n1721;
  wire n1724;
  wire n1727;
  wire n1730;
  wire n1733;
  wire n1736;
  wire n1739;
  wire n1742;
  wire n1745;
  wire n1748;
  wire n1751;
  wire n1754;
  wire n1757;
  wire n1760;
  wire n1763;
  wire n1766;
  wire n1769;
  wire n1772;
  wire n1775;
  wire n1778;
  wire n1781;
  wire n1784;
  wire n1787;
  wire n1790;
  wire n1793;
  wire n1796;
  wire n1799;
  wire n1802;
  wire n1805;
  wire n1808;
  wire n1811;
  wire n1814;
  wire n1817;
  wire n1820;
  wire n1823;
  wire n1826;
  wire n1829;
  wire n1832;
  wire n1835;
  wire n1838;
  wire n1841;
  wire n1844;
  wire n1847;
  wire n1850;
  wire n1853;
  wire n1856;
  wire n1859;
  wire n1862;
  wire n1865;
  wire n1868;
  wire n1871;
  wire n1874;
  wire n1877;
  wire n1880;
  wire n1883;
  wire n1886;
  wire n1889;
  wire n1892;
  wire n1895;
  wire n1898;
  wire n1901;
  wire n1904;
  wire n1907;
  wire n1910;
  wire n1913;
  wire n1916;
  wire n1919;
  wire n1922;
  wire n1925;
  wire n1928;
  wire n1931;
  wire n1934;
  wire n1937;
  wire n1940;
  wire n1943;
  wire n1946;
  wire n1949;
  wire n1952;
  wire n1955;
  wire n1958;
  wire n1961;
  wire n1964;
  wire n1967;
  wire n1970;
  wire n1973;
  wire n1976;
  wire n1979;
  wire n1982;
  wire n1985;
  wire n1988;
  wire n1991;
  wire n1994;
  wire n1997;
  wire n2000;
  wire n2003;
  wire n2006;
  wire n2009;
  wire n2012;
  wire n2015;
  wire n2018;
  wire n2021;
  wire n2024;
  wire n2027;
  wire n2030;
  wire n2033;
  wire n2036;
  wire n2039;
  wire n2042;
  wire n2045;
  wire n2048;
  wire n2051;
  wire n2054;
  wire n2057;
  wire n2060;
  wire n2063;
  wire n2066;
  wire n2069;
  wire n2072;
  wire n2075;
  wire n2078;
  wire n2081;
  wire n2084;
  wire n2087;
  wire n2090;
  wire n2093;
  wire n2096;
  wire n2099;
  wire n2102;
  wire n2105;
  wire n2108;
  wire n2111;
  wire n2114;
  wire n2117;
  wire n2120;
  wire n2123;
  wire n2126;
  wire n2129;
  wire n2132;
  wire n2135;
  wire n2138;
  wire n2141;
  wire n2144;
  wire n2147;
  wire n2150;
  wire n2153;
  wire n2156;
  wire n2159;
  wire n2162;
  wire n2165;
  wire n2168;
  wire n2171;
  wire n2174;
  wire n2177;
  wire n2180;
  wire n2183;
  wire n2186;
  wire n2189;
  wire n2192;
  wire n2195;
  wire n2198;
  wire n2201;
  wire n2204;
  wire n2207;
  wire n2210;
  wire n2213;
  wire n2216;
  wire n2219;
  wire n2222;
  wire n2225;
  wire n2228;
  wire n2231;
  wire n2234;
  wire n2237;
  wire n2240;
  wire n2243;
  wire n2246;
  wire n2249;
  wire n2252;
  wire n2255;
  wire n2258;
  wire n2261;
  wire n2264;
  wire n2267;
  wire n2270;
  wire n2273;
  wire n2276;
  wire n2279;
  wire n2282;
  wire n2285;
  wire n2288;
  wire n2291;
  wire n2294;
  wire [255:0] n2296;
  reg [8:0] n2297;
  assign y = y1; //(module output)
  /* fppowtf32.vhdl:30:8  */
  assign y0 = n2297; // (signal)
  /* fppowtf32.vhdl:32:8  */
  assign y1 = y0; // (signal)
  /* fppowtf32.vhdl:36:19  */
  assign n1529 = x == 8'b00000000;
  /* fppowtf32.vhdl:37:19  */
  assign n1532 = x == 8'b00000001;
  /* fppowtf32.vhdl:38:19  */
  assign n1535 = x == 8'b00000010;
  /* fppowtf32.vhdl:39:19  */
  assign n1538 = x == 8'b00000011;
  /* fppowtf32.vhdl:40:19  */
  assign n1541 = x == 8'b00000100;
  /* fppowtf32.vhdl:41:19  */
  assign n1544 = x == 8'b00000101;
  /* fppowtf32.vhdl:42:19  */
  assign n1547 = x == 8'b00000110;
  /* fppowtf32.vhdl:43:19  */
  assign n1550 = x == 8'b00000111;
  /* fppowtf32.vhdl:44:19  */
  assign n1553 = x == 8'b00001000;
  /* fppowtf32.vhdl:45:19  */
  assign n1556 = x == 8'b00001001;
  /* fppowtf32.vhdl:46:19  */
  assign n1559 = x == 8'b00001010;
  /* fppowtf32.vhdl:47:19  */
  assign n1562 = x == 8'b00001011;
  /* fppowtf32.vhdl:48:19  */
  assign n1565 = x == 8'b00001100;
  /* fppowtf32.vhdl:49:19  */
  assign n1568 = x == 8'b00001101;
  /* fppowtf32.vhdl:50:19  */
  assign n1571 = x == 8'b00001110;
  /* fppowtf32.vhdl:51:19  */
  assign n1574 = x == 8'b00001111;
  /* fppowtf32.vhdl:52:19  */
  assign n1577 = x == 8'b00010000;
  /* fppowtf32.vhdl:53:19  */
  assign n1580 = x == 8'b00010001;
  /* fppowtf32.vhdl:54:19  */
  assign n1583 = x == 8'b00010010;
  /* fppowtf32.vhdl:55:19  */
  assign n1586 = x == 8'b00010011;
  /* fppowtf32.vhdl:56:19  */
  assign n1589 = x == 8'b00010100;
  /* fppowtf32.vhdl:57:19  */
  assign n1592 = x == 8'b00010101;
  /* fppowtf32.vhdl:58:19  */
  assign n1595 = x == 8'b00010110;
  /* fppowtf32.vhdl:59:19  */
  assign n1598 = x == 8'b00010111;
  /* fppowtf32.vhdl:60:19  */
  assign n1601 = x == 8'b00011000;
  /* fppowtf32.vhdl:61:19  */
  assign n1604 = x == 8'b00011001;
  /* fppowtf32.vhdl:62:19  */
  assign n1607 = x == 8'b00011010;
  /* fppowtf32.vhdl:63:19  */
  assign n1610 = x == 8'b00011011;
  /* fppowtf32.vhdl:64:19  */
  assign n1613 = x == 8'b00011100;
  /* fppowtf32.vhdl:65:19  */
  assign n1616 = x == 8'b00011101;
  /* fppowtf32.vhdl:66:19  */
  assign n1619 = x == 8'b00011110;
  /* fppowtf32.vhdl:67:19  */
  assign n1622 = x == 8'b00011111;
  /* fppowtf32.vhdl:68:19  */
  assign n1625 = x == 8'b00100000;
  /* fppowtf32.vhdl:69:19  */
  assign n1628 = x == 8'b00100001;
  /* fppowtf32.vhdl:70:19  */
  assign n1631 = x == 8'b00100010;
  /* fppowtf32.vhdl:71:19  */
  assign n1634 = x == 8'b00100011;
  /* fppowtf32.vhdl:72:19  */
  assign n1637 = x == 8'b00100100;
  /* fppowtf32.vhdl:73:19  */
  assign n1640 = x == 8'b00100101;
  /* fppowtf32.vhdl:74:19  */
  assign n1643 = x == 8'b00100110;
  /* fppowtf32.vhdl:75:19  */
  assign n1646 = x == 8'b00100111;
  /* fppowtf32.vhdl:76:19  */
  assign n1649 = x == 8'b00101000;
  /* fppowtf32.vhdl:77:19  */
  assign n1652 = x == 8'b00101001;
  /* fppowtf32.vhdl:78:19  */
  assign n1655 = x == 8'b00101010;
  /* fppowtf32.vhdl:79:19  */
  assign n1658 = x == 8'b00101011;
  /* fppowtf32.vhdl:80:19  */
  assign n1661 = x == 8'b00101100;
  /* fppowtf32.vhdl:81:19  */
  assign n1664 = x == 8'b00101101;
  /* fppowtf32.vhdl:82:19  */
  assign n1667 = x == 8'b00101110;
  /* fppowtf32.vhdl:83:19  */
  assign n1670 = x == 8'b00101111;
  /* fppowtf32.vhdl:84:19  */
  assign n1673 = x == 8'b00110000;
  /* fppowtf32.vhdl:85:19  */
  assign n1676 = x == 8'b00110001;
  /* fppowtf32.vhdl:86:19  */
  assign n1679 = x == 8'b00110010;
  /* fppowtf32.vhdl:87:19  */
  assign n1682 = x == 8'b00110011;
  /* fppowtf32.vhdl:88:19  */
  assign n1685 = x == 8'b00110100;
  /* fppowtf32.vhdl:89:19  */
  assign n1688 = x == 8'b00110101;
  /* fppowtf32.vhdl:90:19  */
  assign n1691 = x == 8'b00110110;
  /* fppowtf32.vhdl:91:19  */
  assign n1694 = x == 8'b00110111;
  /* fppowtf32.vhdl:92:19  */
  assign n1697 = x == 8'b00111000;
  /* fppowtf32.vhdl:93:19  */
  assign n1700 = x == 8'b00111001;
  /* fppowtf32.vhdl:94:19  */
  assign n1703 = x == 8'b00111010;
  /* fppowtf32.vhdl:95:19  */
  assign n1706 = x == 8'b00111011;
  /* fppowtf32.vhdl:96:19  */
  assign n1709 = x == 8'b00111100;
  /* fppowtf32.vhdl:97:19  */
  assign n1712 = x == 8'b00111101;
  /* fppowtf32.vhdl:98:19  */
  assign n1715 = x == 8'b00111110;
  /* fppowtf32.vhdl:99:19  */
  assign n1718 = x == 8'b00111111;
  /* fppowtf32.vhdl:100:19  */
  assign n1721 = x == 8'b01000000;
  /* fppowtf32.vhdl:101:19  */
  assign n1724 = x == 8'b01000001;
  /* fppowtf32.vhdl:102:19  */
  assign n1727 = x == 8'b01000010;
  /* fppowtf32.vhdl:103:19  */
  assign n1730 = x == 8'b01000011;
  /* fppowtf32.vhdl:104:19  */
  assign n1733 = x == 8'b01000100;
  /* fppowtf32.vhdl:105:19  */
  assign n1736 = x == 8'b01000101;
  /* fppowtf32.vhdl:106:19  */
  assign n1739 = x == 8'b01000110;
  /* fppowtf32.vhdl:107:19  */
  assign n1742 = x == 8'b01000111;
  /* fppowtf32.vhdl:108:19  */
  assign n1745 = x == 8'b01001000;
  /* fppowtf32.vhdl:109:19  */
  assign n1748 = x == 8'b01001001;
  /* fppowtf32.vhdl:110:19  */
  assign n1751 = x == 8'b01001010;
  /* fppowtf32.vhdl:111:19  */
  assign n1754 = x == 8'b01001011;
  /* fppowtf32.vhdl:112:19  */
  assign n1757 = x == 8'b01001100;
  /* fppowtf32.vhdl:113:19  */
  assign n1760 = x == 8'b01001101;
  /* fppowtf32.vhdl:114:19  */
  assign n1763 = x == 8'b01001110;
  /* fppowtf32.vhdl:115:19  */
  assign n1766 = x == 8'b01001111;
  /* fppowtf32.vhdl:116:19  */
  assign n1769 = x == 8'b01010000;
  /* fppowtf32.vhdl:117:19  */
  assign n1772 = x == 8'b01010001;
  /* fppowtf32.vhdl:118:19  */
  assign n1775 = x == 8'b01010010;
  /* fppowtf32.vhdl:119:19  */
  assign n1778 = x == 8'b01010011;
  /* fppowtf32.vhdl:120:19  */
  assign n1781 = x == 8'b01010100;
  /* fppowtf32.vhdl:121:19  */
  assign n1784 = x == 8'b01010101;
  /* fppowtf32.vhdl:122:19  */
  assign n1787 = x == 8'b01010110;
  /* fppowtf32.vhdl:123:19  */
  assign n1790 = x == 8'b01010111;
  /* fppowtf32.vhdl:124:19  */
  assign n1793 = x == 8'b01011000;
  /* fppowtf32.vhdl:125:19  */
  assign n1796 = x == 8'b01011001;
  /* fppowtf32.vhdl:126:19  */
  assign n1799 = x == 8'b01011010;
  /* fppowtf32.vhdl:127:19  */
  assign n1802 = x == 8'b01011011;
  /* fppowtf32.vhdl:128:19  */
  assign n1805 = x == 8'b01011100;
  /* fppowtf32.vhdl:129:19  */
  assign n1808 = x == 8'b01011101;
  /* fppowtf32.vhdl:130:19  */
  assign n1811 = x == 8'b01011110;
  /* fppowtf32.vhdl:131:19  */
  assign n1814 = x == 8'b01011111;
  /* fppowtf32.vhdl:132:19  */
  assign n1817 = x == 8'b01100000;
  /* fppowtf32.vhdl:133:19  */
  assign n1820 = x == 8'b01100001;
  /* fppowtf32.vhdl:134:19  */
  assign n1823 = x == 8'b01100010;
  /* fppowtf32.vhdl:135:19  */
  assign n1826 = x == 8'b01100011;
  /* fppowtf32.vhdl:136:19  */
  assign n1829 = x == 8'b01100100;
  /* fppowtf32.vhdl:137:19  */
  assign n1832 = x == 8'b01100101;
  /* fppowtf32.vhdl:138:19  */
  assign n1835 = x == 8'b01100110;
  /* fppowtf32.vhdl:139:19  */
  assign n1838 = x == 8'b01100111;
  /* fppowtf32.vhdl:140:19  */
  assign n1841 = x == 8'b01101000;
  /* fppowtf32.vhdl:141:19  */
  assign n1844 = x == 8'b01101001;
  /* fppowtf32.vhdl:142:19  */
  assign n1847 = x == 8'b01101010;
  /* fppowtf32.vhdl:143:19  */
  assign n1850 = x == 8'b01101011;
  /* fppowtf32.vhdl:144:19  */
  assign n1853 = x == 8'b01101100;
  /* fppowtf32.vhdl:145:19  */
  assign n1856 = x == 8'b01101101;
  /* fppowtf32.vhdl:146:19  */
  assign n1859 = x == 8'b01101110;
  /* fppowtf32.vhdl:147:19  */
  assign n1862 = x == 8'b01101111;
  /* fppowtf32.vhdl:148:19  */
  assign n1865 = x == 8'b01110000;
  /* fppowtf32.vhdl:149:19  */
  assign n1868 = x == 8'b01110001;
  /* fppowtf32.vhdl:150:19  */
  assign n1871 = x == 8'b01110010;
  /* fppowtf32.vhdl:151:19  */
  assign n1874 = x == 8'b01110011;
  /* fppowtf32.vhdl:152:19  */
  assign n1877 = x == 8'b01110100;
  /* fppowtf32.vhdl:153:19  */
  assign n1880 = x == 8'b01110101;
  /* fppowtf32.vhdl:154:19  */
  assign n1883 = x == 8'b01110110;
  /* fppowtf32.vhdl:155:19  */
  assign n1886 = x == 8'b01110111;
  /* fppowtf32.vhdl:156:19  */
  assign n1889 = x == 8'b01111000;
  /* fppowtf32.vhdl:157:19  */
  assign n1892 = x == 8'b01111001;
  /* fppowtf32.vhdl:158:19  */
  assign n1895 = x == 8'b01111010;
  /* fppowtf32.vhdl:159:19  */
  assign n1898 = x == 8'b01111011;
  /* fppowtf32.vhdl:160:19  */
  assign n1901 = x == 8'b01111100;
  /* fppowtf32.vhdl:161:19  */
  assign n1904 = x == 8'b01111101;
  /* fppowtf32.vhdl:162:19  */
  assign n1907 = x == 8'b01111110;
  /* fppowtf32.vhdl:163:19  */
  assign n1910 = x == 8'b01111111;
  /* fppowtf32.vhdl:164:19  */
  assign n1913 = x == 8'b10000000;
  /* fppowtf32.vhdl:165:19  */
  assign n1916 = x == 8'b10000001;
  /* fppowtf32.vhdl:166:19  */
  assign n1919 = x == 8'b10000010;
  /* fppowtf32.vhdl:167:19  */
  assign n1922 = x == 8'b10000011;
  /* fppowtf32.vhdl:168:19  */
  assign n1925 = x == 8'b10000100;
  /* fppowtf32.vhdl:169:19  */
  assign n1928 = x == 8'b10000101;
  /* fppowtf32.vhdl:170:19  */
  assign n1931 = x == 8'b10000110;
  /* fppowtf32.vhdl:171:19  */
  assign n1934 = x == 8'b10000111;
  /* fppowtf32.vhdl:172:19  */
  assign n1937 = x == 8'b10001000;
  /* fppowtf32.vhdl:173:19  */
  assign n1940 = x == 8'b10001001;
  /* fppowtf32.vhdl:174:19  */
  assign n1943 = x == 8'b10001010;
  /* fppowtf32.vhdl:175:19  */
  assign n1946 = x == 8'b10001011;
  /* fppowtf32.vhdl:176:19  */
  assign n1949 = x == 8'b10001100;
  /* fppowtf32.vhdl:177:19  */
  assign n1952 = x == 8'b10001101;
  /* fppowtf32.vhdl:178:19  */
  assign n1955 = x == 8'b10001110;
  /* fppowtf32.vhdl:179:19  */
  assign n1958 = x == 8'b10001111;
  /* fppowtf32.vhdl:180:19  */
  assign n1961 = x == 8'b10010000;
  /* fppowtf32.vhdl:181:19  */
  assign n1964 = x == 8'b10010001;
  /* fppowtf32.vhdl:182:19  */
  assign n1967 = x == 8'b10010010;
  /* fppowtf32.vhdl:183:19  */
  assign n1970 = x == 8'b10010011;
  /* fppowtf32.vhdl:184:19  */
  assign n1973 = x == 8'b10010100;
  /* fppowtf32.vhdl:185:19  */
  assign n1976 = x == 8'b10010101;
  /* fppowtf32.vhdl:186:19  */
  assign n1979 = x == 8'b10010110;
  /* fppowtf32.vhdl:187:19  */
  assign n1982 = x == 8'b10010111;
  /* fppowtf32.vhdl:188:19  */
  assign n1985 = x == 8'b10011000;
  /* fppowtf32.vhdl:189:19  */
  assign n1988 = x == 8'b10011001;
  /* fppowtf32.vhdl:190:19  */
  assign n1991 = x == 8'b10011010;
  /* fppowtf32.vhdl:191:19  */
  assign n1994 = x == 8'b10011011;
  /* fppowtf32.vhdl:192:19  */
  assign n1997 = x == 8'b10011100;
  /* fppowtf32.vhdl:193:19  */
  assign n2000 = x == 8'b10011101;
  /* fppowtf32.vhdl:194:19  */
  assign n2003 = x == 8'b10011110;
  /* fppowtf32.vhdl:195:19  */
  assign n2006 = x == 8'b10011111;
  /* fppowtf32.vhdl:196:19  */
  assign n2009 = x == 8'b10100000;
  /* fppowtf32.vhdl:197:19  */
  assign n2012 = x == 8'b10100001;
  /* fppowtf32.vhdl:198:19  */
  assign n2015 = x == 8'b10100010;
  /* fppowtf32.vhdl:199:19  */
  assign n2018 = x == 8'b10100011;
  /* fppowtf32.vhdl:200:19  */
  assign n2021 = x == 8'b10100100;
  /* fppowtf32.vhdl:201:19  */
  assign n2024 = x == 8'b10100101;
  /* fppowtf32.vhdl:202:19  */
  assign n2027 = x == 8'b10100110;
  /* fppowtf32.vhdl:203:19  */
  assign n2030 = x == 8'b10100111;
  /* fppowtf32.vhdl:204:19  */
  assign n2033 = x == 8'b10101000;
  /* fppowtf32.vhdl:205:19  */
  assign n2036 = x == 8'b10101001;
  /* fppowtf32.vhdl:206:19  */
  assign n2039 = x == 8'b10101010;
  /* fppowtf32.vhdl:207:19  */
  assign n2042 = x == 8'b10101011;
  /* fppowtf32.vhdl:208:19  */
  assign n2045 = x == 8'b10101100;
  /* fppowtf32.vhdl:209:19  */
  assign n2048 = x == 8'b10101101;
  /* fppowtf32.vhdl:210:19  */
  assign n2051 = x == 8'b10101110;
  /* fppowtf32.vhdl:211:19  */
  assign n2054 = x == 8'b10101111;
  /* fppowtf32.vhdl:212:19  */
  assign n2057 = x == 8'b10110000;
  /* fppowtf32.vhdl:213:19  */
  assign n2060 = x == 8'b10110001;
  /* fppowtf32.vhdl:214:19  */
  assign n2063 = x == 8'b10110010;
  /* fppowtf32.vhdl:215:19  */
  assign n2066 = x == 8'b10110011;
  /* fppowtf32.vhdl:216:19  */
  assign n2069 = x == 8'b10110100;
  /* fppowtf32.vhdl:217:19  */
  assign n2072 = x == 8'b10110101;
  /* fppowtf32.vhdl:218:19  */
  assign n2075 = x == 8'b10110110;
  /* fppowtf32.vhdl:219:19  */
  assign n2078 = x == 8'b10110111;
  /* fppowtf32.vhdl:220:19  */
  assign n2081 = x == 8'b10111000;
  /* fppowtf32.vhdl:221:19  */
  assign n2084 = x == 8'b10111001;
  /* fppowtf32.vhdl:222:19  */
  assign n2087 = x == 8'b10111010;
  /* fppowtf32.vhdl:223:19  */
  assign n2090 = x == 8'b10111011;
  /* fppowtf32.vhdl:224:19  */
  assign n2093 = x == 8'b10111100;
  /* fppowtf32.vhdl:225:19  */
  assign n2096 = x == 8'b10111101;
  /* fppowtf32.vhdl:226:19  */
  assign n2099 = x == 8'b10111110;
  /* fppowtf32.vhdl:227:19  */
  assign n2102 = x == 8'b10111111;
  /* fppowtf32.vhdl:228:19  */
  assign n2105 = x == 8'b11000000;
  /* fppowtf32.vhdl:229:19  */
  assign n2108 = x == 8'b11000001;
  /* fppowtf32.vhdl:230:19  */
  assign n2111 = x == 8'b11000010;
  /* fppowtf32.vhdl:231:19  */
  assign n2114 = x == 8'b11000011;
  /* fppowtf32.vhdl:232:19  */
  assign n2117 = x == 8'b11000100;
  /* fppowtf32.vhdl:233:19  */
  assign n2120 = x == 8'b11000101;
  /* fppowtf32.vhdl:234:19  */
  assign n2123 = x == 8'b11000110;
  /* fppowtf32.vhdl:235:19  */
  assign n2126 = x == 8'b11000111;
  /* fppowtf32.vhdl:236:19  */
  assign n2129 = x == 8'b11001000;
  /* fppowtf32.vhdl:237:19  */
  assign n2132 = x == 8'b11001001;
  /* fppowtf32.vhdl:238:19  */
  assign n2135 = x == 8'b11001010;
  /* fppowtf32.vhdl:239:19  */
  assign n2138 = x == 8'b11001011;
  /* fppowtf32.vhdl:240:19  */
  assign n2141 = x == 8'b11001100;
  /* fppowtf32.vhdl:241:19  */
  assign n2144 = x == 8'b11001101;
  /* fppowtf32.vhdl:242:19  */
  assign n2147 = x == 8'b11001110;
  /* fppowtf32.vhdl:243:19  */
  assign n2150 = x == 8'b11001111;
  /* fppowtf32.vhdl:244:19  */
  assign n2153 = x == 8'b11010000;
  /* fppowtf32.vhdl:245:19  */
  assign n2156 = x == 8'b11010001;
  /* fppowtf32.vhdl:246:19  */
  assign n2159 = x == 8'b11010010;
  /* fppowtf32.vhdl:247:19  */
  assign n2162 = x == 8'b11010011;
  /* fppowtf32.vhdl:248:19  */
  assign n2165 = x == 8'b11010100;
  /* fppowtf32.vhdl:249:19  */
  assign n2168 = x == 8'b11010101;
  /* fppowtf32.vhdl:250:19  */
  assign n2171 = x == 8'b11010110;
  /* fppowtf32.vhdl:251:19  */
  assign n2174 = x == 8'b11010111;
  /* fppowtf32.vhdl:252:19  */
  assign n2177 = x == 8'b11011000;
  /* fppowtf32.vhdl:253:19  */
  assign n2180 = x == 8'b11011001;
  /* fppowtf32.vhdl:254:19  */
  assign n2183 = x == 8'b11011010;
  /* fppowtf32.vhdl:255:19  */
  assign n2186 = x == 8'b11011011;
  /* fppowtf32.vhdl:256:19  */
  assign n2189 = x == 8'b11011100;
  /* fppowtf32.vhdl:257:19  */
  assign n2192 = x == 8'b11011101;
  /* fppowtf32.vhdl:258:19  */
  assign n2195 = x == 8'b11011110;
  /* fppowtf32.vhdl:259:19  */
  assign n2198 = x == 8'b11011111;
  /* fppowtf32.vhdl:260:19  */
  assign n2201 = x == 8'b11100000;
  /* fppowtf32.vhdl:261:19  */
  assign n2204 = x == 8'b11100001;
  /* fppowtf32.vhdl:262:19  */
  assign n2207 = x == 8'b11100010;
  /* fppowtf32.vhdl:263:19  */
  assign n2210 = x == 8'b11100011;
  /* fppowtf32.vhdl:264:19  */
  assign n2213 = x == 8'b11100100;
  /* fppowtf32.vhdl:265:19  */
  assign n2216 = x == 8'b11100101;
  /* fppowtf32.vhdl:266:19  */
  assign n2219 = x == 8'b11100110;
  /* fppowtf32.vhdl:267:19  */
  assign n2222 = x == 8'b11100111;
  /* fppowtf32.vhdl:268:19  */
  assign n2225 = x == 8'b11101000;
  /* fppowtf32.vhdl:269:19  */
  assign n2228 = x == 8'b11101001;
  /* fppowtf32.vhdl:270:19  */
  assign n2231 = x == 8'b11101010;
  /* fppowtf32.vhdl:271:19  */
  assign n2234 = x == 8'b11101011;
  /* fppowtf32.vhdl:272:19  */
  assign n2237 = x == 8'b11101100;
  /* fppowtf32.vhdl:273:19  */
  assign n2240 = x == 8'b11101101;
  /* fppowtf32.vhdl:274:19  */
  assign n2243 = x == 8'b11101110;
  /* fppowtf32.vhdl:275:19  */
  assign n2246 = x == 8'b11101111;
  /* fppowtf32.vhdl:276:19  */
  assign n2249 = x == 8'b11110000;
  /* fppowtf32.vhdl:277:19  */
  assign n2252 = x == 8'b11110001;
  /* fppowtf32.vhdl:278:19  */
  assign n2255 = x == 8'b11110010;
  /* fppowtf32.vhdl:279:19  */
  assign n2258 = x == 8'b11110011;
  /* fppowtf32.vhdl:280:19  */
  assign n2261 = x == 8'b11110100;
  /* fppowtf32.vhdl:281:19  */
  assign n2264 = x == 8'b11110101;
  /* fppowtf32.vhdl:282:19  */
  assign n2267 = x == 8'b11110110;
  /* fppowtf32.vhdl:283:19  */
  assign n2270 = x == 8'b11110111;
  /* fppowtf32.vhdl:284:19  */
  assign n2273 = x == 8'b11111000;
  /* fppowtf32.vhdl:285:19  */
  assign n2276 = x == 8'b11111001;
  /* fppowtf32.vhdl:286:19  */
  assign n2279 = x == 8'b11111010;
  /* fppowtf32.vhdl:287:19  */
  assign n2282 = x == 8'b11111011;
  /* fppowtf32.vhdl:288:19  */
  assign n2285 = x == 8'b11111100;
  /* fppowtf32.vhdl:289:19  */
  assign n2288 = x == 8'b11111101;
  /* fppowtf32.vhdl:290:19  */
  assign n2291 = x == 8'b11111110;
  /* fppowtf32.vhdl:291:19  */
  assign n2294 = x == 8'b11111111;
  assign n2296 = {n2294, n2291, n2288, n2285, n2282, n2279, n2276, n2273, n2270, n2267, n2264, n2261, n2258, n2255, n2252, n2249, n2246, n2243, n2240, n2237, n2234, n2231, n2228, n2225, n2222, n2219, n2216, n2213, n2210, n2207, n2204, n2201, n2198, n2195, n2192, n2189, n2186, n2183, n2180, n2177, n2174, n2171, n2168, n2165, n2162, n2159, n2156, n2153, n2150, n2147, n2144, n2141, n2138, n2135, n2132, n2129, n2126, n2123, n2120, n2117, n2114, n2111, n2108, n2105, n2102, n2099, n2096, n2093, n2090, n2087, n2084, n2081, n2078, n2075, n2072, n2069, n2066, n2063, n2060, n2057, n2054, n2051, n2048, n2045, n2042, n2039, n2036, n2033, n2030, n2027, n2024, n2021, n2018, n2015, n2012, n2009, n2006, n2003, n2000, n1997, n1994, n1991, n1988, n1985, n1982, n1979, n1976, n1973, n1970, n1967, n1964, n1961, n1958, n1955, n1952, n1949, n1946, n1943, n1940, n1937, n1934, n1931, n1928, n1925, n1922, n1919, n1916, n1913, n1910, n1907, n1904, n1901, n1898, n1895, n1892, n1889, n1886, n1883, n1880, n1877, n1874, n1871, n1868, n1865, n1862, n1859, n1856, n1853, n1850, n1847, n1844, n1841, n1838, n1835, n1832, n1829, n1826, n1823, n1820, n1817, n1814, n1811, n1808, n1805, n1802, n1799, n1796, n1793, n1790, n1787, n1784, n1781, n1778, n1775, n1772, n1769, n1766, n1763, n1760, n1757, n1754, n1751, n1748, n1745, n1742, n1739, n1736, n1733, n1730, n1727, n1724, n1721, n1718, n1715, n1712, n1709, n1706, n1703, n1700, n1697, n1694, n1691, n1688, n1685, n1682, n1679, n1676, n1673, n1670, n1667, n1664, n1661, n1658, n1655, n1652, n1649, n1646, n1643, n1640, n1637, n1634, n1631, n1628, n1625, n1622, n1619, n1616, n1613, n1610, n1607, n1604, n1601, n1598, n1595, n1592, n1589, n1586, n1583, n1580, n1577, n1574, n1571, n1568, n1565, n1562, n1559, n1556, n1553, n1550, n1547, n1544, n1541, n1538, n1535, n1532, n1529};
  /* fppowtf32.vhdl:35:4  */
  always @*
    case (n2296)
      256'b1000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2297 = 9'b100000001;
      256'b0100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2297 = 9'b100000010;
      256'b0010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2297 = 9'b100000010;
      256'b0001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2297 = 9'b100000011;
      256'b0000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2297 = 9'b100000011;
      256'b0000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2297 = 9'b100000100;
      256'b0000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2297 = 9'b100000100;
      256'b0000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2297 = 9'b100000101;
      256'b0000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2297 = 9'b100000101;
      256'b0000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2297 = 9'b100000110;
      256'b0000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2297 = 9'b100000110;
      256'b0000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2297 = 9'b100000111;
      256'b0000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2297 = 9'b100000111;
      256'b0000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2297 = 9'b100001000;
      256'b0000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2297 = 9'b100001000;
      256'b0000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2297 = 9'b100001001;
      256'b0000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2297 = 9'b100001001;
      256'b0000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2297 = 9'b100001010;
      256'b0000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2297 = 9'b100001010;
      256'b0000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2297 = 9'b100001011;
      256'b0000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2297 = 9'b100001011;
      256'b0000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2297 = 9'b100001100;
      256'b0000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2297 = 9'b100001101;
      256'b0000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2297 = 9'b100001101;
      256'b0000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2297 = 9'b100001110;
      256'b0000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2297 = 9'b100001110;
      256'b0000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2297 = 9'b100001111;
      256'b0000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2297 = 9'b100001111;
      256'b0000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2297 = 9'b100010000;
      256'b0000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2297 = 9'b100010000;
      256'b0000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2297 = 9'b100010001;
      256'b0000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2297 = 9'b100010010;
      256'b0000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2297 = 9'b100010010;
      256'b0000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2297 = 9'b100010011;
      256'b0000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2297 = 9'b100010011;
      256'b0000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2297 = 9'b100010100;
      256'b0000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2297 = 9'b100010100;
      256'b0000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2297 = 9'b100010101;
      256'b0000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2297 = 9'b100010110;
      256'b0000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2297 = 9'b100010110;
      256'b0000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2297 = 9'b100010111;
      256'b0000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2297 = 9'b100010111;
      256'b0000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2297 = 9'b100011000;
      256'b0000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2297 = 9'b100011001;
      256'b0000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2297 = 9'b100011001;
      256'b0000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2297 = 9'b100011010;
      256'b0000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2297 = 9'b100011010;
      256'b0000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2297 = 9'b100011011;
      256'b0000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2297 = 9'b100011100;
      256'b0000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2297 = 9'b100011100;
      256'b0000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2297 = 9'b100011101;
      256'b0000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2297 = 9'b100011101;
      256'b0000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2297 = 9'b100011110;
      256'b0000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2297 = 9'b100011111;
      256'b0000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2297 = 9'b100011111;
      256'b0000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2297 = 9'b100100000;
      256'b0000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2297 = 9'b100100001;
      256'b0000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2297 = 9'b100100001;
      256'b0000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2297 = 9'b100100010;
      256'b0000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2297 = 9'b100100010;
      256'b0000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2297 = 9'b100100011;
      256'b0000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2297 = 9'b100100100;
      256'b0000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2297 = 9'b100100100;
      256'b0000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2297 = 9'b100100101;
      256'b0000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2297 = 9'b100100110;
      256'b0000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2297 = 9'b100100110;
      256'b0000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2297 = 9'b100100111;
      256'b0000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2297 = 9'b100101000;
      256'b0000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2297 = 9'b100101000;
      256'b0000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2297 = 9'b100101001;
      256'b0000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2297 = 9'b100101010;
      256'b0000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2297 = 9'b100101010;
      256'b0000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2297 = 9'b100101011;
      256'b0000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2297 = 9'b100101100;
      256'b0000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2297 = 9'b100101100;
      256'b0000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2297 = 9'b100101101;
      256'b0000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2297 = 9'b100101110;
      256'b0000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2297 = 9'b100101111;
      256'b0000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2297 = 9'b100101111;
      256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2297 = 9'b100110000;
      256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2297 = 9'b100110001;
      256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2297 = 9'b100110001;
      256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2297 = 9'b100110010;
      256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2297 = 9'b100110011;
      256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2297 = 9'b100110011;
      256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2297 = 9'b100110100;
      256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2297 = 9'b100110101;
      256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2297 = 9'b100110110;
      256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2297 = 9'b100110110;
      256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2297 = 9'b100110111;
      256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2297 = 9'b100111000;
      256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2297 = 9'b100111001;
      256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2297 = 9'b100111001;
      256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2297 = 9'b100111010;
      256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2297 = 9'b100111011;
      256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2297 = 9'b100111100;
      256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2297 = 9'b100111100;
      256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2297 = 9'b100111101;
      256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2297 = 9'b100111110;
      256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2297 = 9'b100111111;
      256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2297 = 9'b100111111;
      256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2297 = 9'b101000000;
      256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2297 = 9'b101000001;
      256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2297 = 9'b101000010;
      256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2297 = 9'b101000011;
      256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2297 = 9'b101000011;
      256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2297 = 9'b101000100;
      256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2297 = 9'b101000101;
      256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2297 = 9'b101000110;
      256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2297 = 9'b101000111;
      256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2297 = 9'b101000111;
      256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2297 = 9'b101001000;
      256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2297 = 9'b101001001;
      256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2297 = 9'b101001010;
      256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2297 = 9'b101001011;
      256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2297 = 9'b101001011;
      256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2297 = 9'b101001100;
      256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2297 = 9'b101001101;
      256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2297 = 9'b101001110;
      256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2297 = 9'b101001111;
      256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2297 = 9'b101010000;
      256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2297 = 9'b101010001;
      256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2297 = 9'b101010001;
      256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2297 = 9'b101010010;
      256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2297 = 9'b101010011;
      256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2297 = 9'b101010100;
      256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2297 = 9'b101010101;
      256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2297 = 9'b101010110;
      256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2297 = 9'b010101100;
      256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2297 = 9'b010101100;
      256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2297 = 9'b010101101;
      256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2297 = 9'b010101101;
      256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2297 = 9'b010101101;
      256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2297 = 9'b010101110;
      256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2297 = 9'b010101110;
      256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2297 = 9'b010101111;
      256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2297 = 9'b010101111;
      256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2297 = 9'b010110000;
      256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2297 = 9'b010110000;
      256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2297 = 9'b010110001;
      256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2297 = 9'b010110001;
      256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2297 = 9'b010110010;
      256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2297 = 9'b010110010;
      256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2297 = 9'b010110011;
      256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2297 = 9'b010110011;
      256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2297 = 9'b010110100;
      256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2297 = 9'b010110100;
      256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2297 = 9'b010110101;
      256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2297 = 9'b010110101;
      256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2297 = 9'b010110110;
      256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2297 = 9'b010110110;
      256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2297 = 9'b010110111;
      256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2297 = 9'b010110111;
      256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2297 = 9'b010111000;
      256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2297 = 9'b010111000;
      256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2297 = 9'b010111001;
      256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2297 = 9'b010111001;
      256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2297 = 9'b010111010;
      256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2297 = 9'b010111010;
      256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2297 = 9'b010111011;
      256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2297 = 9'b010111011;
      256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2297 = 9'b010111100;
      256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2297 = 9'b010111100;
      256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2297 = 9'b010111101;
      256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2297 = 9'b010111101;
      256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2297 = 9'b010111110;
      256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2297 = 9'b010111110;
      256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2297 = 9'b010111111;
      256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2297 = 9'b011000000;
      256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2297 = 9'b011000000;
      256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2297 = 9'b011000001;
      256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2297 = 9'b011000001;
      256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2297 = 9'b011000010;
      256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2297 = 9'b011000010;
      256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000: n2297 = 9'b011000011;
      256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000: n2297 = 9'b011000100;
      256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000: n2297 = 9'b011000100;
      256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000: n2297 = 9'b011000101;
      256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000: n2297 = 9'b011000101;
      256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000: n2297 = 9'b011000110;
      256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000: n2297 = 9'b011000110;
      256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000: n2297 = 9'b011000111;
      256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000: n2297 = 9'b011001000;
      256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000: n2297 = 9'b011001000;
      256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000: n2297 = 9'b011001001;
      256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000: n2297 = 9'b011001010;
      256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000: n2297 = 9'b011001010;
      256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000: n2297 = 9'b011001011;
      256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000: n2297 = 9'b011001011;
      256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000: n2297 = 9'b011001100;
      256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000: n2297 = 9'b011001101;
      256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000: n2297 = 9'b011001101;
      256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000: n2297 = 9'b011001110;
      256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000: n2297 = 9'b011001111;
      256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000: n2297 = 9'b011001111;
      256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000: n2297 = 9'b011010000;
      256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000: n2297 = 9'b011010001;
      256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000: n2297 = 9'b011010001;
      256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000: n2297 = 9'b011010010;
      256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000: n2297 = 9'b011010011;
      256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000: n2297 = 9'b011010011;
      256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000: n2297 = 9'b011010100;
      256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000: n2297 = 9'b011010101;
      256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000: n2297 = 9'b011010101;
      256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000: n2297 = 9'b011010110;
      256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000: n2297 = 9'b011010111;
      256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000: n2297 = 9'b011010111;
      256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000: n2297 = 9'b011011000;
      256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000: n2297 = 9'b011011001;
      256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000: n2297 = 9'b011011010;
      256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000: n2297 = 9'b011011010;
      256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000: n2297 = 9'b011011011;
      256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000: n2297 = 9'b011011100;
      256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000: n2297 = 9'b011011100;
      256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000: n2297 = 9'b011011101;
      256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000: n2297 = 9'b011011110;
      256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000: n2297 = 9'b011011111;
      256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000: n2297 = 9'b011011111;
      256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000: n2297 = 9'b011100000;
      256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000: n2297 = 9'b011100001;
      256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000: n2297 = 9'b011100010;
      256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000: n2297 = 9'b011100010;
      256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000: n2297 = 9'b011100011;
      256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000: n2297 = 9'b011100100;
      256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000: n2297 = 9'b011100101;
      256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000: n2297 = 9'b011100110;
      256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000: n2297 = 9'b011100110;
      256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000: n2297 = 9'b011100111;
      256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000: n2297 = 9'b011101000;
      256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000: n2297 = 9'b011101001;
      256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000: n2297 = 9'b011101010;
      256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000: n2297 = 9'b011101011;
      256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000: n2297 = 9'b011101011;
      256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000: n2297 = 9'b011101100;
      256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000: n2297 = 9'b011101101;
      256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000: n2297 = 9'b011101110;
      256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000: n2297 = 9'b011101111;
      256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000: n2297 = 9'b011110000;
      256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000: n2297 = 9'b011110001;
      256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000: n2297 = 9'b011110001;
      256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000: n2297 = 9'b011110010;
      256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000: n2297 = 9'b011110011;
      256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000: n2297 = 9'b011110100;
      256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000: n2297 = 9'b011110101;
      256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000: n2297 = 9'b011110110;
      256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000: n2297 = 9'b011110111;
      256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000: n2297 = 9'b011111000;
      256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000: n2297 = 9'b011111001;
      256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000: n2297 = 9'b011111010;
      256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000: n2297 = 9'b011111011;
      256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000: n2297 = 9'b011111100;
      256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000: n2297 = 9'b011111101;
      256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000: n2297 = 9'b011111110;
      256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100: n2297 = 9'b011111111;
      256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010: n2297 = 9'b100000000;
      256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001: n2297 = 9'b100000000;
      default: n2297 = 9'bX;
    endcase
endmodule

module leftshifter11_by_max_11_freq500_uid13
  (input  clk,
   input  [10:0] x,
   input  [3:0] s,
   output [21:0] r);
  wire [3:0] ps;
  wire [3:0] ps_d1;
  wire [10:0] level0;
  wire [10:0] level0_d1;
  wire [10:0] level0_d2;
  wire [10:0] level0_d3;
  wire [11:0] level1;
  wire [11:0] level1_d1;
  wire [13:0] level2;
  wire [17:0] level3;
  wire [25:0] level4;
  wire [11:0] n1497;
  wire n1498;
  wire [11:0] n1499;
  wire [11:0] n1501;
  wire [13:0] n1503;
  wire n1504;
  wire [13:0] n1505;
  wire [13:0] n1507;
  wire [17:0] n1509;
  wire n1510;
  wire [17:0] n1511;
  wire [17:0] n1513;
  wire [25:0] n1515;
  wire n1516;
  wire [25:0] n1517;
  wire [25:0] n1519;
  wire [21:0] n1520;
  reg [3:0] n1521;
  reg [10:0] n1522;
  reg [10:0] n1523;
  reg [10:0] n1524;
  reg [11:0] n1525;
  assign r = n1520; //(module output)
  /* fppowtf32.vhdl:2433:12  */
  assign ps_d1 = n1521; // (signal)
  /* fppowtf32.vhdl:2435:16  */
  assign level0_d1 = n1522; // (signal)
  /* fppowtf32.vhdl:2435:27  */
  assign level0_d2 = n1523; // (signal)
  /* fppowtf32.vhdl:2435:38  */
  assign level0_d3 = n1524; // (signal)
  /* fppowtf32.vhdl:2437:8  */
  assign level1 = n1499; // (signal)
  /* fppowtf32.vhdl:2437:16  */
  assign level1_d1 = n1525; // (signal)
  /* fppowtf32.vhdl:2439:8  */
  assign level2 = n1505; // (signal)
  /* fppowtf32.vhdl:2441:8  */
  assign level3 = n1511; // (signal)
  /* fppowtf32.vhdl:2443:8  */
  assign level4 = n1517; // (signal)
  /* fppowtf32.vhdl:2458:23  */
  assign n1497 = {level0_d3, 1'b0};
  /* fppowtf32.vhdl:2458:52  */
  assign n1498 = ps[0]; // extract
  /* fppowtf32.vhdl:2458:45  */
  assign n1499 = n1498 ? n1497 : n1501;
  /* fppowtf32.vhdl:2458:90  */
  assign n1501 = {1'b0, level0_d3};
  /* fppowtf32.vhdl:2459:23  */
  assign n1503 = {level1_d1, 2'b00};
  /* fppowtf32.vhdl:2459:55  */
  assign n1504 = ps_d1[1]; // extract
  /* fppowtf32.vhdl:2459:45  */
  assign n1505 = n1504 ? n1503 : n1507;
  /* fppowtf32.vhdl:2459:93  */
  assign n1507 = {2'b00, level1_d1};
  /* fppowtf32.vhdl:2460:20  */
  assign n1509 = {level2, 4'b0000};
  /* fppowtf32.vhdl:2460:52  */
  assign n1510 = ps_d1[2]; // extract
  /* fppowtf32.vhdl:2460:42  */
  assign n1511 = n1510 ? n1509 : n1513;
  /* fppowtf32.vhdl:2460:90  */
  assign n1513 = {4'b0000, level2};
  /* fppowtf32.vhdl:2461:20  */
  assign n1515 = {level3, 8'b00000000};
  /* fppowtf32.vhdl:2461:52  */
  assign n1516 = ps_d1[3]; // extract
  /* fppowtf32.vhdl:2461:42  */
  assign n1517 = n1516 ? n1515 : n1519;
  /* fppowtf32.vhdl:2461:90  */
  assign n1519 = {8'b00000000, level3};
  /* fppowtf32.vhdl:2462:15  */
  assign n1520 = level4[21:0]; // extract
  /* fppowtf32.vhdl:2448:10  */
  always @(posedge clk)
    n1521 <= ps;
  /* fppowtf32.vhdl:2448:10  */
  always @(posedge clk)
    n1522 <= level0;
  /* fppowtf32.vhdl:2448:10  */
  always @(posedge clk)
    n1523 <= level0_d1;
  /* fppowtf32.vhdl:2448:10  */
  always @(posedge clk)
    n1524 <= level0_d2;
  /* fppowtf32.vhdl:2448:10  */
  always @(posedge clk)
    n1525 <= level1;
endmodule

module lzoc_20_freq500_uid11
  (input  clk,
   input  [19:0] i,
   input  ozb,
   output [4:0] o);
  wire sozb;
  wire sozb_d1;
  wire sozb_d2;
  wire [30:0] level5;
  wire [30:0] level5_d1;
  wire digit4;
  wire digit4_d1;
  wire digit4_d2;
  wire [14:0] level4;
  wire [14:0] level4_d1;
  wire digit3;
  wire digit3_d1;
  wire [6:0] level3;
  wire digit2;
  wire [2:0] level2;
  wire [2:0] level2_d1;
  wire [2:0] z;
  wire [1:0] lowbits;
  wire [2:0] outhighbits;
  wire [2:0] outhighbits_d1;
  wire ozb_d1;
  wire ozb_d2;
  wire ozb_d3;
  wire n1403;
  wire n1404;
  wire n1405;
  wire n1406;
  wire n1407;
  wire n1408;
  wire n1409;
  wire n1410;
  wire n1411;
  wire n1412;
  wire n1413;
  wire [3:0] n1414;
  wire [3:0] n1415;
  wire [2:0] n1416;
  wire [10:0] n1417;
  wire [30:0] n1418;
  wire [15:0] n1420;
  wire [3:0] n1421;
  wire [3:0] n1422;
  wire [3:0] n1423;
  wire [3:0] n1424;
  wire [15:0] n1425;
  wire n1426;
  wire n1427;
  wire [14:0] n1429;
  wire [14:0] n1430;
  wire [14:0] n1431;
  wire [7:0] n1433;
  wire [3:0] n1434;
  wire [3:0] n1435;
  wire [7:0] n1436;
  wire n1437;
  wire n1438;
  wire [6:0] n1440;
  wire [6:0] n1441;
  wire [6:0] n1442;
  wire [3:0] n1444;
  wire [3:0] n1445;
  wire n1446;
  wire n1447;
  wire [2:0] n1449;
  wire [2:0] n1450;
  wire [2:0] n1451;
  wire n1452;
  wire [2:0] n1453;
  wire [2:0] n1454;
  wire n1457;
  wire n1460;
  wire n1463;
  wire n1466;
  wire [3:0] n1468;
  reg [1:0] n1469;
  wire [1:0] n1470;
  wire [2:0] n1471;
  wire [4:0] n1473;
  reg n1474;
  reg n1475;
  reg [30:0] n1476;
  reg n1477;
  reg n1478;
  reg [14:0] n1479;
  reg n1480;
  reg [2:0] n1481;
  reg [2:0] n1482;
  reg n1483;
  reg n1484;
  reg n1485;
  assign o = n1473; //(module output)
  /* fppowtf32.vhdl:2338:8  */
  assign sozb = ozb; // (signal)
  /* fppowtf32.vhdl:2338:14  */
  assign sozb_d1 = n1474; // (signal)
  /* fppowtf32.vhdl:2338:23  */
  assign sozb_d2 = n1475; // (signal)
  /* fppowtf32.vhdl:2340:8  */
  assign level5 = n1418; // (signal)
  /* fppowtf32.vhdl:2340:16  */
  assign level5_d1 = n1476; // (signal)
  /* fppowtf32.vhdl:2342:8  */
  assign digit4 = n1427; // (signal)
  /* fppowtf32.vhdl:2342:16  */
  assign digit4_d1 = n1477; // (signal)
  /* fppowtf32.vhdl:2342:27  */
  assign digit4_d2 = n1478; // (signal)
  /* fppowtf32.vhdl:2344:8  */
  assign level4 = n1430; // (signal)
  /* fppowtf32.vhdl:2344:16  */
  assign level4_d1 = n1479; // (signal)
  /* fppowtf32.vhdl:2346:8  */
  assign digit3 = n1438; // (signal)
  /* fppowtf32.vhdl:2346:16  */
  assign digit3_d1 = n1480; // (signal)
  /* fppowtf32.vhdl:2348:8  */
  assign level3 = n1441; // (signal)
  /* fppowtf32.vhdl:2350:8  */
  assign digit2 = n1447; // (signal)
  /* fppowtf32.vhdl:2352:8  */
  assign level2 = n1450; // (signal)
  /* fppowtf32.vhdl:2352:16  */
  assign level2_d1 = n1481; // (signal)
  /* fppowtf32.vhdl:2354:8  */
  assign z = n1453; // (signal)
  /* fppowtf32.vhdl:2356:8  */
  assign lowbits = n1469; // (signal)
  /* fppowtf32.vhdl:2358:8  */
  assign outhighbits = n1471; // (signal)
  /* fppowtf32.vhdl:2358:21  */
  assign outhighbits_d1 = n1482; // (signal)
  /* fppowtf32.vhdl:2360:8  */
  assign ozb_d1 = n1483; // (signal)
  /* fppowtf32.vhdl:2360:16  */
  assign ozb_d2 = n1484; // (signal)
  /* fppowtf32.vhdl:2360:24  */
  assign ozb_d3 = n1485; // (signal)
  /* fppowtf32.vhdl:2382:34  */
  assign n1403 = ~sozb;
  /* fppowtf32.vhdl:2382:34  */
  assign n1404 = ~sozb;
  /* fppowtf32.vhdl:2382:34  */
  assign n1405 = ~sozb;
  /* fppowtf32.vhdl:2382:34  */
  assign n1406 = ~sozb;
  /* fppowtf32.vhdl:2382:34  */
  assign n1407 = ~sozb;
  /* fppowtf32.vhdl:2382:34  */
  assign n1408 = ~sozb;
  /* fppowtf32.vhdl:2382:34  */
  assign n1409 = ~sozb;
  /* fppowtf32.vhdl:2382:34  */
  assign n1410 = ~sozb;
  /* fppowtf32.vhdl:2382:34  */
  assign n1411 = ~sozb;
  /* fppowtf32.vhdl:2382:34  */
  assign n1412 = ~sozb;
  /* fppowtf32.vhdl:2382:34  */
  assign n1413 = ~sozb;
  assign n1414 = {n1413, n1412, n1411, n1410};
  assign n1415 = {n1409, n1408, n1407, n1406};
  assign n1416 = {n1405, n1404, n1403};
  assign n1417 = {n1414, n1415, n1416};
  /* fppowtf32.vhdl:2382:16  */
  assign n1418 = {i, n1417};
  /* fppowtf32.vhdl:2384:28  */
  assign n1420 = level5[30:15]; // extract
  assign n1421 = {sozb, sozb, sozb, sozb};
  assign n1422 = {sozb, sozb, sozb, sozb};
  assign n1423 = {sozb, sozb, sozb, sozb};
  assign n1424 = {sozb, sozb, sozb, sozb};
  assign n1425 = {n1421, n1422, n1423, n1424};
  /* fppowtf32.vhdl:2384:43  */
  assign n1426 = n1420 == n1425;
  /* fppowtf32.vhdl:2384:17  */
  assign n1427 = n1426 ? 1'b1 : 1'b0;
  /* fppowtf32.vhdl:2385:22  */
  assign n1429 = level5_d1[14:0]; // extract
  /* fppowtf32.vhdl:2385:36  */
  assign n1430 = digit4_d1 ? n1429 : n1431;
  /* fppowtf32.vhdl:2385:69  */
  assign n1431 = level5_d1[30:16]; // extract
  /* fppowtf32.vhdl:2386:28  */
  assign n1433 = level4[14:7]; // extract
  assign n1434 = {sozb_d1, sozb_d1, sozb_d1, sozb_d1};
  assign n1435 = {sozb_d1, sozb_d1, sozb_d1, sozb_d1};
  assign n1436 = {n1434, n1435};
  /* fppowtf32.vhdl:2386:42  */
  assign n1437 = n1433 == n1436;
  /* fppowtf32.vhdl:2386:17  */
  assign n1438 = n1437 ? 1'b1 : 1'b0;
  /* fppowtf32.vhdl:2387:22  */
  assign n1440 = level4_d1[6:0]; // extract
  /* fppowtf32.vhdl:2387:35  */
  assign n1441 = digit3_d1 ? n1440 : n1442;
  /* fppowtf32.vhdl:2387:68  */
  assign n1442 = level4_d1[14:8]; // extract
  /* fppowtf32.vhdl:2388:28  */
  assign n1444 = level3[6:3]; // extract
  assign n1445 = {sozb_d2, sozb_d2, sozb_d2, sozb_d2};
  /* fppowtf32.vhdl:2388:41  */
  assign n1446 = n1444 == n1445;
  /* fppowtf32.vhdl:2388:17  */
  assign n1447 = n1446 ? 1'b1 : 1'b0;
  /* fppowtf32.vhdl:2389:19  */
  assign n1449 = level3[2:0]; // extract
  /* fppowtf32.vhdl:2389:32  */
  assign n1450 = digit2 ? n1449 : n1451;
  /* fppowtf32.vhdl:2389:59  */
  assign n1451 = level3[6:4]; // extract
  /* fppowtf32.vhdl:2391:30  */
  assign n1452 = ~ozb_d3;
  /* fppowtf32.vhdl:2391:19  */
  assign n1453 = n1452 ? level2_d1 : n1454;
  /* fppowtf32.vhdl:2391:41  */
  assign n1454 = ~level2_d1;
  /* fppowtf32.vhdl:2393:12  */
  assign n1457 = z == 3'b000;
  /* fppowtf32.vhdl:2394:12  */
  assign n1460 = z == 3'b001;
  /* fppowtf32.vhdl:2395:12  */
  assign n1463 = z == 3'b010;
  /* fppowtf32.vhdl:2396:12  */
  assign n1466 = z == 3'b011;
  assign n1468 = {n1466, n1463, n1460, n1457};
  /* fppowtf32.vhdl:2392:4  */
  always @*
    case (n1468)
      4'b1000: n1469 = 2'b01;
      4'b0100: n1469 = 2'b01;
      4'b0010: n1469 = 2'b10;
      4'b0001: n1469 = 2'b11;
      default: n1469 = 2'b00;
    endcase
  /* fppowtf32.vhdl:2398:29  */
  assign n1470 = {digit4_d2, digit3_d1};
  /* fppowtf32.vhdl:2398:50  */
  assign n1471 = {n1470, digit2};
  /* fppowtf32.vhdl:2399:24  */
  assign n1473 = {outhighbits_d1, lowbits};
  /* fppowtf32.vhdl:2365:10  */
  always @(posedge clk)
    n1474 <= sozb;
  /* fppowtf32.vhdl:2365:10  */
  always @(posedge clk)
    n1475 <= sozb_d1;
  /* fppowtf32.vhdl:2365:10  */
  always @(posedge clk)
    n1476 <= level5;
  /* fppowtf32.vhdl:2365:10  */
  always @(posedge clk)
    n1477 <= digit4;
  /* fppowtf32.vhdl:2365:10  */
  always @(posedge clk)
    n1478 <= digit4_d1;
  /* fppowtf32.vhdl:2365:10  */
  always @(posedge clk)
    n1479 <= level4;
  /* fppowtf32.vhdl:2365:10  */
  always @(posedge clk)
    n1480 <= digit3;
  /* fppowtf32.vhdl:2365:10  */
  always @(posedge clk)
    n1481 <= level2;
  /* fppowtf32.vhdl:2365:10  */
  always @(posedge clk)
    n1482 <= outhighbits;
  /* fppowtf32.vhdl:2365:10  */
  always @(posedge clk)
    n1483 <= ozb;
  /* fppowtf32.vhdl:2365:10  */
  always @(posedge clk)
    n1484 <= ozb_d1;
  /* fppowtf32.vhdl:2365:10  */
  always @(posedge clk)
    n1485 <= ozb_d2;
endmodule

module fpexp_8_10_freq500_uid71
  (input  clk,
   input  [31:0] x,
   output [20:0] r);
  wire [1:0] xexn;
  wire [1:0] xexn_d1;
  wire [1:0] xexn_d2;
  wire [1:0] xexn_d3;
  wire [1:0] xexn_d4;
  wire [1:0] xexn_d5;
  wire [1:0] xexn_d6;
  wire [1:0] xexn_d7;
  wire xsign;
  wire xsign_d1;
  wire xsign_d2;
  wire xsign_d3;
  wire xsign_d4;
  wire xsign_d5;
  wire xsign_d6;
  wire xsign_d7;
  wire [7:0] xexpfield;
  wire [7:0] xexpfield_d1;
  wire [20:0] xfrac;
  wire [9:0] e0;
  wire [9:0] e0_d1;
  wire [9:0] e0_d2;
  wire [9:0] e0_d3;
  wire [9:0] e0_d4;
  wire [9:0] e0_d5;
  wire [9:0] e0_d6;
  wire [9:0] e0_d7;
  wire [9:0] e0_d8;
  wire [9:0] e0_d9;
  wire [9:0] e0_d10;
  wire [9:0] e0_d11;
  wire [9:0] e0_d12;
  wire [9:0] e0_d13;
  wire [9:0] e0_d14;
  wire [9:0] shiftval;
  wire [9:0] shiftval_d1;
  wire resultwillbeone;
  wire resultwillbeone_d1;
  wire [21:0] mxu;
  wire [8:0] maxshift;
  wire [8:0] maxshift_d1;
  wire [8:0] maxshift_d2;
  wire [8:0] maxshift_d3;
  wire [8:0] maxshift_d4;
  wire [8:0] maxshift_d5;
  wire [8:0] maxshift_d6;
  wire [8:0] maxshift_d7;
  wire [8:0] maxshift_d8;
  wire [8:0] maxshift_d9;
  wire [8:0] maxshift_d10;
  wire [8:0] maxshift_d11;
  wire [8:0] maxshift_d12;
  wire [8:0] maxshift_d13;
  wire [8:0] maxshift_d14;
  wire [8:0] maxshift_d15;
  wire overflow0;
  wire [4:0] shiftvalin;
  wire [40:0] fixx0;
  wire [19:0] ufixx;
  wire [13:0] expy;
  wire [8:0] k;
  wire [8:0] k_d1;
  wire [8:0] k_d2;
  wire neednonorm;
  wire [19:0] preroundbiassig;
  wire roundbit;
  wire [19:0] roundnormaddend;
  wire [19:0] roundedexpsigres;
  wire [19:0] roundedexpsig;
  wire ofl1;
  wire ofl1_d1;
  wire ofl1_d2;
  wire ofl1_d3;
  wire ofl1_d4;
  wire ofl1_d5;
  wire ofl2;
  wire ofl3;
  wire ofl3_d1;
  wire ofl3_d2;
  wire ofl3_d3;
  wire ofl3_d4;
  wire ofl3_d5;
  wire ofl3_d6;
  wire ofl3_d7;
  wire ofl;
  wire ufl1;
  wire ufl2;
  wire ufl2_d1;
  wire ufl2_d2;
  wire ufl2_d3;
  wire ufl2_d4;
  wire ufl2_d5;
  wire ufl2_d6;
  wire ufl2_d7;
  wire ufl3;
  wire ufl3_d1;
  wire ufl3_d2;
  wire ufl3_d3;
  wire ufl3_d4;
  wire ufl3_d5;
  wire ufl;
  wire [1:0] rexn;
  wire [1:0] n1198;
  wire n1199;
  wire [7:0] n1200;
  wire [20:0] n1201;
  wire [9:0] n1204;
  wire [9:0] n1205;
  wire n1206;
  wire [21:0] n1208;
  wire n1210;
  wire n1211;
  wire [8:0] n1212;
  wire n1213;
  wire n1214;
  wire [4:0] n1216;
  wire [40:0] mantissa_shift_n1217;
  wire [19:0] n1220;
  wire n1221;
  wire [19:0] n1222;
  wire [13:0] exp_helper_n1224;
  wire [8:0] exp_helper_n1225;
  wire n1230;
  wire [9:0] n1231;
  wire [19:0] n1233;
  wire [19:0] n1234;
  wire [9:0] n1235;
  wire [19:0] n1237;
  wire n1238;
  wire n1239;
  wire n1240;
  wire n1241;
  wire [9:0] n1242;
  wire [18:0] n1244;
  wire [19:0] n1245;
  localparam n1246 = 1'b0;
  wire [19:0] roundedexpsigoperandadder_n1247;
  wire n1251;
  wire [19:0] n1252;
  wire n1254;
  wire n1255;
  wire n1256;
  wire n1257;
  wire n1258;
  wire n1259;
  wire n1260;
  wire n1261;
  wire n1262;
  wire n1263;
  wire n1264;
  wire n1265;
  wire n1266;
  wire n1267;
  wire n1268;
  wire n1269;
  wire n1270;
  wire n1271;
  wire n1272;
  wire n1273;
  wire n1274;
  wire n1275;
  wire n1276;
  wire n1277;
  wire n1278;
  wire n1279;
  wire n1280;
  wire n1281;
  wire n1282;
  wire n1283;
  wire n1284;
  wire n1285;
  wire n1286;
  wire n1287;
  wire n1288;
  wire n1289;
  wire n1290;
  wire n1291;
  wire n1292;
  wire n1293;
  wire n1294;
  wire n1295;
  wire n1296;
  wire n1297;
  wire n1298;
  wire n1299;
  wire n1300;
  wire n1303;
  wire [1:0] n1304;
  wire [1:0] n1306;
  wire [1:0] n1308;
  wire [2:0] n1311;
  wire [17:0] n1312;
  wire [20:0] n1313;
  reg [1:0] n1314;
  reg [1:0] n1315;
  reg [1:0] n1316;
  reg [1:0] n1317;
  reg [1:0] n1318;
  reg [1:0] n1319;
  reg [1:0] n1320;
  reg n1321;
  reg n1322;
  reg n1323;
  reg n1324;
  reg n1325;
  reg n1326;
  reg n1327;
  reg [7:0] n1328;
  reg [9:0] n1329;
  reg [9:0] n1330;
  reg [9:0] n1331;
  reg [9:0] n1332;
  reg [9:0] n1333;
  reg [9:0] n1334;
  reg [9:0] n1335;
  reg [9:0] n1336;
  reg [9:0] n1337;
  reg [9:0] n1338;
  reg [9:0] n1339;
  reg [9:0] n1340;
  reg [9:0] n1341;
  reg [9:0] n1342;
  reg [9:0] n1343;
  reg n1344;
  reg [8:0] n1345;
  reg [8:0] n1346;
  reg [8:0] n1347;
  reg [8:0] n1348;
  reg [8:0] n1349;
  reg [8:0] n1350;
  reg [8:0] n1351;
  reg [8:0] n1352;
  reg [8:0] n1353;
  reg [8:0] n1354;
  reg [8:0] n1355;
  reg [8:0] n1356;
  reg [8:0] n1357;
  reg [8:0] n1358;
  reg [8:0] n1359;
  reg [8:0] n1360;
  reg [8:0] n1361;
  reg n1362;
  reg n1363;
  reg n1364;
  reg n1365;
  reg n1366;
  reg n1367;
  reg n1368;
  reg n1369;
  reg n1370;
  reg n1371;
  reg n1372;
  reg n1373;
  reg n1374;
  reg n1375;
  reg n1376;
  reg n1377;
  reg n1378;
  reg n1379;
  reg n1380;
  reg n1381;
  reg n1382;
  reg n1383;
  reg n1384;
  reg n1385;
  assign r = n1313; //(module output)
  /* fppowtf32.vhdl:5529:8  */
  assign xexn = n1198; // (signal)
  /* fppowtf32.vhdl:5529:14  */
  assign xexn_d1 = n1314; // (signal)
  /* fppowtf32.vhdl:5529:23  */
  assign xexn_d2 = n1315; // (signal)
  /* fppowtf32.vhdl:5529:32  */
  assign xexn_d3 = n1316; // (signal)
  /* fppowtf32.vhdl:5529:41  */
  assign xexn_d4 = n1317; // (signal)
  /* fppowtf32.vhdl:5529:50  */
  assign xexn_d5 = n1318; // (signal)
  /* fppowtf32.vhdl:5529:59  */
  assign xexn_d6 = n1319; // (signal)
  /* fppowtf32.vhdl:5529:68  */
  assign xexn_d7 = n1320; // (signal)
  /* fppowtf32.vhdl:5531:8  */
  assign xsign = n1199; // (signal)
  /* fppowtf32.vhdl:5531:15  */
  assign xsign_d1 = n1321; // (signal)
  /* fppowtf32.vhdl:5531:25  */
  assign xsign_d2 = n1322; // (signal)
  /* fppowtf32.vhdl:5531:35  */
  assign xsign_d3 = n1323; // (signal)
  /* fppowtf32.vhdl:5531:45  */
  assign xsign_d4 = n1324; // (signal)
  /* fppowtf32.vhdl:5531:55  */
  assign xsign_d5 = n1325; // (signal)
  /* fppowtf32.vhdl:5531:65  */
  assign xsign_d6 = n1326; // (signal)
  /* fppowtf32.vhdl:5531:75  */
  assign xsign_d7 = n1327; // (signal)
  /* fppowtf32.vhdl:5533:8  */
  assign xexpfield = n1200; // (signal)
  /* fppowtf32.vhdl:5533:19  */
  assign xexpfield_d1 = n1328; // (signal)
  /* fppowtf32.vhdl:5535:8  */
  assign xfrac = n1201; // (signal)
  /* fppowtf32.vhdl:5537:8  */
  assign e0 = 10'b0001110010; // (signal)
  /* fppowtf32.vhdl:5537:12  */
  assign e0_d1 = n1329; // (signal)
  /* fppowtf32.vhdl:5537:19  */
  assign e0_d2 = n1330; // (signal)
  /* fppowtf32.vhdl:5537:26  */
  assign e0_d3 = n1331; // (signal)
  /* fppowtf32.vhdl:5537:33  */
  assign e0_d4 = n1332; // (signal)
  /* fppowtf32.vhdl:5537:40  */
  assign e0_d5 = n1333; // (signal)
  /* fppowtf32.vhdl:5537:47  */
  assign e0_d6 = n1334; // (signal)
  /* fppowtf32.vhdl:5537:54  */
  assign e0_d7 = n1335; // (signal)
  /* fppowtf32.vhdl:5537:61  */
  assign e0_d8 = n1336; // (signal)
  /* fppowtf32.vhdl:5537:68  */
  assign e0_d9 = n1337; // (signal)
  /* fppowtf32.vhdl:5537:75  */
  assign e0_d10 = n1338; // (signal)
  /* fppowtf32.vhdl:5537:83  */
  assign e0_d11 = n1339; // (signal)
  /* fppowtf32.vhdl:5537:91  */
  assign e0_d12 = n1340; // (signal)
  /* fppowtf32.vhdl:5537:99  */
  assign e0_d13 = n1341; // (signal)
  /* fppowtf32.vhdl:5537:107  */
  assign e0_d14 = n1342; // (signal)
  /* fppowtf32.vhdl:5539:8  */
  assign shiftval = n1205; // (signal)
  /* fppowtf32.vhdl:5539:18  */
  assign shiftval_d1 = n1343; // (signal)
  /* fppowtf32.vhdl:5541:8  */
  assign resultwillbeone = n1206; // (signal)
  /* fppowtf32.vhdl:5541:25  */
  assign resultwillbeone_d1 = n1344; // (signal)
  /* fppowtf32.vhdl:5543:8  */
  assign mxu = n1208; // (signal)
  /* fppowtf32.vhdl:5545:8  */
  assign maxshift = 9'b000010011; // (signal)
  /* fppowtf32.vhdl:5545:18  */
  assign maxshift_d1 = n1345; // (signal)
  /* fppowtf32.vhdl:5545:31  */
  assign maxshift_d2 = n1346; // (signal)
  /* fppowtf32.vhdl:5545:44  */
  assign maxshift_d3 = n1347; // (signal)
  /* fppowtf32.vhdl:5545:57  */
  assign maxshift_d4 = n1348; // (signal)
  /* fppowtf32.vhdl:5545:70  */
  assign maxshift_d5 = n1349; // (signal)
  /* fppowtf32.vhdl:5545:83  */
  assign maxshift_d6 = n1350; // (signal)
  /* fppowtf32.vhdl:5545:96  */
  assign maxshift_d7 = n1351; // (signal)
  /* fppowtf32.vhdl:5545:109  */
  assign maxshift_d8 = n1352; // (signal)
  /* fppowtf32.vhdl:5545:122  */
  assign maxshift_d9 = n1353; // (signal)
  /* fppowtf32.vhdl:5545:135  */
  assign maxshift_d10 = n1354; // (signal)
  /* fppowtf32.vhdl:5545:149  */
  assign maxshift_d11 = n1355; // (signal)
  /* fppowtf32.vhdl:5545:163  */
  assign maxshift_d12 = n1356; // (signal)
  /* fppowtf32.vhdl:5545:177  */
  assign maxshift_d13 = n1357; // (signal)
  /* fppowtf32.vhdl:5545:191  */
  assign maxshift_d14 = n1358; // (signal)
  /* fppowtf32.vhdl:5545:205  */
  assign maxshift_d15 = n1359; // (signal)
  /* fppowtf32.vhdl:5547:8  */
  assign overflow0 = n1214; // (signal)
  /* fppowtf32.vhdl:5549:8  */
  assign shiftvalin = n1216; // (signal)
  /* fppowtf32.vhdl:5551:8  */
  assign fixx0 = mantissa_shift_n1217; // (signal)
  /* fppowtf32.vhdl:5553:8  */
  assign ufixx = n1222; // (signal)
  /* fppowtf32.vhdl:5555:8  */
  assign expy = exp_helper_n1224; // (signal)
  /* fppowtf32.vhdl:5557:8  */
  assign k = exp_helper_n1225; // (signal)
  /* fppowtf32.vhdl:5557:11  */
  assign k_d1 = n1360; // (signal)
  /* fppowtf32.vhdl:5557:17  */
  assign k_d2 = n1361; // (signal)
  /* fppowtf32.vhdl:5559:8  */
  assign neednonorm = n1230; // (signal)
  /* fppowtf32.vhdl:5561:8  */
  assign preroundbiassig = n1234; // (signal)
  /* fppowtf32.vhdl:5563:8  */
  assign roundbit = n1239; // (signal)
  /* fppowtf32.vhdl:5565:8  */
  assign roundnormaddend = n1245; // (signal)
  /* fppowtf32.vhdl:5567:8  */
  assign roundedexpsigres = roundedexpsigoperandadder_n1247; // (signal)
  /* fppowtf32.vhdl:5569:8  */
  assign roundedexpsig = n1252; // (signal)
  /* fppowtf32.vhdl:5571:8  */
  assign ofl1 = n1260; // (signal)
  /* fppowtf32.vhdl:5571:14  */
  assign ofl1_d1 = n1362; // (signal)
  /* fppowtf32.vhdl:5571:23  */
  assign ofl1_d2 = n1363; // (signal)
  /* fppowtf32.vhdl:5571:32  */
  assign ofl1_d3 = n1364; // (signal)
  /* fppowtf32.vhdl:5571:41  */
  assign ofl1_d4 = n1365; // (signal)
  /* fppowtf32.vhdl:5571:50  */
  assign ofl1_d5 = n1366; // (signal)
  /* fppowtf32.vhdl:5573:8  */
  assign ofl2 = n1271; // (signal)
  /* fppowtf32.vhdl:5575:8  */
  assign ofl3 = n1277; // (signal)
  /* fppowtf32.vhdl:5575:14  */
  assign ofl3_d1 = n1367; // (signal)
  /* fppowtf32.vhdl:5575:23  */
  assign ofl3_d2 = n1368; // (signal)
  /* fppowtf32.vhdl:5575:32  */
  assign ofl3_d3 = n1369; // (signal)
  /* fppowtf32.vhdl:5575:41  */
  assign ofl3_d4 = n1370; // (signal)
  /* fppowtf32.vhdl:5575:50  */
  assign ofl3_d5 = n1371; // (signal)
  /* fppowtf32.vhdl:5575:59  */
  assign ofl3_d6 = n1372; // (signal)
  /* fppowtf32.vhdl:5575:68  */
  assign ofl3_d7 = n1373; // (signal)
  /* fppowtf32.vhdl:5577:8  */
  assign ofl = n1279; // (signal)
  /* fppowtf32.vhdl:5579:8  */
  assign ufl1 = n1287; // (signal)
  /* fppowtf32.vhdl:5581:8  */
  assign ufl2 = n1292; // (signal)
  /* fppowtf32.vhdl:5581:14  */
  assign ufl2_d1 = n1374; // (signal)
  /* fppowtf32.vhdl:5581:23  */
  assign ufl2_d2 = n1375; // (signal)
  /* fppowtf32.vhdl:5581:32  */
  assign ufl2_d3 = n1376; // (signal)
  /* fppowtf32.vhdl:5581:41  */
  assign ufl2_d4 = n1377; // (signal)
  /* fppowtf32.vhdl:5581:50  */
  assign ufl2_d5 = n1378; // (signal)
  /* fppowtf32.vhdl:5581:59  */
  assign ufl2_d6 = n1379; // (signal)
  /* fppowtf32.vhdl:5581:68  */
  assign ufl2_d7 = n1380; // (signal)
  /* fppowtf32.vhdl:5583:8  */
  assign ufl3 = n1298; // (signal)
  /* fppowtf32.vhdl:5583:14  */
  assign ufl3_d1 = n1381; // (signal)
  /* fppowtf32.vhdl:5583:23  */
  assign ufl3_d2 = n1382; // (signal)
  /* fppowtf32.vhdl:5583:32  */
  assign ufl3_d3 = n1383; // (signal)
  /* fppowtf32.vhdl:5583:41  */
  assign ufl3_d4 = n1384; // (signal)
  /* fppowtf32.vhdl:5583:50  */
  assign ufl3_d5 = n1385; // (signal)
  /* fppowtf32.vhdl:5585:8  */
  assign ufl = n1300; // (signal)
  /* fppowtf32.vhdl:5587:8  */
  assign rexn = n1304; // (signal)
  /* fppowtf32.vhdl:5671:13  */
  assign n1198 = x[31:30]; // extract
  /* fppowtf32.vhdl:5672:14  */
  assign n1199 = x[29]; // extract
  /* fppowtf32.vhdl:5673:18  */
  assign n1200 = x[28:21]; // extract
  /* fppowtf32.vhdl:5674:23  */
  assign n1201 = x[20:0]; // extract
  /* fppowtf32.vhdl:5676:22  */
  assign n1204 = {2'b00, xexpfield_d1};
  /* fppowtf32.vhdl:5676:38  */
  assign n1205 = n1204 - e0_d14;
  /* fppowtf32.vhdl:5678:31  */
  assign n1206 = shiftval[9]; // extract
  /* fppowtf32.vhdl:5680:15  */
  assign n1208 = {1'b1, xfrac};
  /* fppowtf32.vhdl:5683:32  */
  assign n1210 = shiftval_d1[9]; // extract
  /* fppowtf32.vhdl:5683:17  */
  assign n1211 = ~n1210;
  /* fppowtf32.vhdl:5683:55  */
  assign n1212 = shiftval_d1[8:0]; // extract
  /* fppowtf32.vhdl:5683:69  */
  assign n1213 = $unsigned(n1212) > $unsigned(maxshift_d15);
  /* fppowtf32.vhdl:5683:39  */
  assign n1214 = n1213 ? n1211 : 1'b0;
  /* fppowtf32.vhdl:5684:26  */
  assign n1216 = shiftval[4:0]; // extract
  /* fppowtf32.vhdl:5685:4  */
  leftshifter22_by_max_19_freq500_uid73 mantissa_shift (
    .clk(clk),
    .x(mxu),
    .s(shiftvalin),
    .r(mantissa_shift_n1217));
  /* fppowtf32.vhdl:5690:28  */
  assign n1220 = fixx0[40:21]; // extract
  /* fppowtf32.vhdl:5690:67  */
  assign n1221 = ~resultwillbeone_d1;
  /* fppowtf32.vhdl:5690:44  */
  assign n1222 = n1221 ? n1220 : 20'b00000000000000000000;
  /* fppowtf32.vhdl:5691:4  */
  exp_8_10_freq500_uid75 exp_helper (
    .clk(clk),
    .ufixx_i(ufixx),
    .xsign(xsign),
    .expy(exp_helper_n1224),
    .k(exp_helper_n1225));
  /* fppowtf32.vhdl:5697:22  */
  assign n1230 = expy[13]; // extract
  /* fppowtf32.vhdl:5699:63  */
  assign n1231 = expy[12:3]; // extract
  /* fppowtf32.vhdl:5699:57  */
  assign n1233 = {10'b0001111111, n1231};
  /* fppowtf32.vhdl:5699:77  */
  assign n1234 = neednonorm ? n1233 : n1237;
  /* fppowtf32.vhdl:5700:52  */
  assign n1235 = expy[11:2]; // extract
  /* fppowtf32.vhdl:5700:46  */
  assign n1237 = {10'b0001111110, n1235};
  /* fppowtf32.vhdl:5701:20  */
  assign n1238 = expy[2]; // extract
  /* fppowtf32.vhdl:5701:25  */
  assign n1239 = neednonorm ? n1238 : n1240;
  /* fppowtf32.vhdl:5701:59  */
  assign n1240 = expy[1]; // extract
  /* fppowtf32.vhdl:5702:27  */
  assign n1241 = k_d2[8]; // extract
  /* fppowtf32.vhdl:5702:31  */
  assign n1242 = {n1241, k_d2};
  /* fppowtf32.vhdl:5702:38  */
  assign n1244 = {n1242, 9'b000000000};
  /* fppowtf32.vhdl:5702:60  */
  assign n1245 = {n1244, roundbit};
  /* fppowtf32.vhdl:5703:4  */
  intadder_20_freq500_uid121 roundedexpsigoperandadder (
    .clk(clk),
    .x(preroundbiassig),
    .y(roundnormaddend),
    .cin(n1246),
    .r(roundedexpsigoperandadder_n1247));
  /* fppowtf32.vhdl:5709:50  */
  assign n1251 = xexn_d7 == 2'b01;
  /* fppowtf32.vhdl:5709:38  */
  assign n1252 = n1251 ? roundedexpsigres : 20'b00011111110000000000;
  /* fppowtf32.vhdl:5710:12  */
  assign n1254 = ~xsign_d2;
  /* fppowtf32.vhdl:5710:25  */
  assign n1255 = n1254 & overflow0;
  /* fppowtf32.vhdl:5710:55  */
  assign n1256 = xexn_d2[1]; // extract
  /* fppowtf32.vhdl:5710:44  */
  assign n1257 = ~n1256;
  /* fppowtf32.vhdl:5710:70  */
  assign n1258 = xexn_d2[0]; // extract
  /* fppowtf32.vhdl:5710:59  */
  assign n1259 = n1257 & n1258;
  /* fppowtf32.vhdl:5710:39  */
  assign n1260 = n1255 & n1259;
  /* fppowtf32.vhdl:5711:12  */
  assign n1261 = ~xsign_d7;
  /* fppowtf32.vhdl:5711:43  */
  assign n1262 = roundedexpsig[18]; // extract
  /* fppowtf32.vhdl:5711:72  */
  assign n1263 = roundedexpsig[19]; // extract
  /* fppowtf32.vhdl:5711:55  */
  assign n1264 = ~n1263;
  /* fppowtf32.vhdl:5711:51  */
  assign n1265 = n1262 & n1264;
  /* fppowtf32.vhdl:5711:25  */
  assign n1266 = n1261 & n1265;
  /* fppowtf32.vhdl:5711:99  */
  assign n1267 = xexn_d7[1]; // extract
  /* fppowtf32.vhdl:5711:88  */
  assign n1268 = ~n1267;
  /* fppowtf32.vhdl:5711:114  */
  assign n1269 = xexn_d7[0]; // extract
  /* fppowtf32.vhdl:5711:103  */
  assign n1270 = n1268 & n1269;
  /* fppowtf32.vhdl:5711:83  */
  assign n1271 = n1266 & n1270;
  /* fppowtf32.vhdl:5712:12  */
  assign n1272 = ~xsign;
  /* fppowtf32.vhdl:5712:30  */
  assign n1273 = xexn[1]; // extract
  /* fppowtf32.vhdl:5712:22  */
  assign n1274 = n1272 & n1273;
  /* fppowtf32.vhdl:5712:46  */
  assign n1275 = xexn[0]; // extract
  /* fppowtf32.vhdl:5712:38  */
  assign n1276 = ~n1275;
  /* fppowtf32.vhdl:5712:34  */
  assign n1277 = n1274 & n1276;
  /* fppowtf32.vhdl:5713:19  */
  assign n1278 = ofl1_d5 | ofl2;
  /* fppowtf32.vhdl:5713:27  */
  assign n1279 = n1278 | ofl3_d7;
  /* fppowtf32.vhdl:5714:26  */
  assign n1280 = roundedexpsig[18]; // extract
  /* fppowtf32.vhdl:5714:51  */
  assign n1281 = roundedexpsig[19]; // extract
  /* fppowtf32.vhdl:5714:34  */
  assign n1282 = n1280 & n1281;
  /* fppowtf32.vhdl:5714:79  */
  assign n1283 = xexn_d7[1]; // extract
  /* fppowtf32.vhdl:5714:68  */
  assign n1284 = ~n1283;
  /* fppowtf32.vhdl:5714:94  */
  assign n1285 = xexn_d7[0]; // extract
  /* fppowtf32.vhdl:5714:83  */
  assign n1286 = n1284 & n1285;
  /* fppowtf32.vhdl:5714:63  */
  assign n1287 = n1282 & n1286;
  /* fppowtf32.vhdl:5715:26  */
  assign n1288 = xexn[1]; // extract
  /* fppowtf32.vhdl:5715:18  */
  assign n1289 = xsign & n1288;
  /* fppowtf32.vhdl:5715:42  */
  assign n1290 = xexn[0]; // extract
  /* fppowtf32.vhdl:5715:34  */
  assign n1291 = ~n1290;
  /* fppowtf32.vhdl:5715:30  */
  assign n1292 = n1289 & n1291;
  /* fppowtf32.vhdl:5716:21  */
  assign n1293 = xsign_d2 & overflow0;
  /* fppowtf32.vhdl:5716:52  */
  assign n1294 = xexn_d2[1]; // extract
  /* fppowtf32.vhdl:5716:41  */
  assign n1295 = ~n1294;
  /* fppowtf32.vhdl:5716:67  */
  assign n1296 = xexn_d2[0]; // extract
  /* fppowtf32.vhdl:5716:56  */
  assign n1297 = n1295 & n1296;
  /* fppowtf32.vhdl:5716:36  */
  assign n1298 = n1293 & n1297;
  /* fppowtf32.vhdl:5717:16  */
  assign n1299 = ufl1 | ufl2_d7;
  /* fppowtf32.vhdl:5717:27  */
  assign n1300 = n1299 | ufl3_d5;
  /* fppowtf32.vhdl:5718:30  */
  assign n1303 = xexn_d7 == 2'b11;
  /* fppowtf32.vhdl:5718:17  */
  assign n1304 = n1303 ? 2'b11 : n1306;
  /* fppowtf32.vhdl:5719:7  */
  assign n1306 = ofl ? 2'b10 : n1308;
  /* fppowtf32.vhdl:5720:7  */
  assign n1308 = ufl ? 2'b00 : 2'b01;
  /* fppowtf32.vhdl:5722:14  */
  assign n1311 = {rexn, 1'b0};
  /* fppowtf32.vhdl:5722:35  */
  assign n1312 = roundedexpsig[17:0]; // extract
  /* fppowtf32.vhdl:5722:20  */
  assign n1313 = {n1311, n1312};
  /* fppowtf32.vhdl:5596:10  */
  always @(posedge clk)
    n1314 <= xexn;
  /* fppowtf32.vhdl:5596:10  */
  always @(posedge clk)
    n1315 <= xexn_d1;
  /* fppowtf32.vhdl:5596:10  */
  always @(posedge clk)
    n1316 <= xexn_d2;
  /* fppowtf32.vhdl:5596:10  */
  always @(posedge clk)
    n1317 <= xexn_d3;
  /* fppowtf32.vhdl:5596:10  */
  always @(posedge clk)
    n1318 <= xexn_d4;
  /* fppowtf32.vhdl:5596:10  */
  always @(posedge clk)
    n1319 <= xexn_d5;
  /* fppowtf32.vhdl:5596:10  */
  always @(posedge clk)
    n1320 <= xexn_d6;
  /* fppowtf32.vhdl:5596:10  */
  always @(posedge clk)
    n1321 <= xsign;
  /* fppowtf32.vhdl:5596:10  */
  always @(posedge clk)
    n1322 <= xsign_d1;
  /* fppowtf32.vhdl:5596:10  */
  always @(posedge clk)
    n1323 <= xsign_d2;
  /* fppowtf32.vhdl:5596:10  */
  always @(posedge clk)
    n1324 <= xsign_d3;
  /* fppowtf32.vhdl:5596:10  */
  always @(posedge clk)
    n1325 <= xsign_d4;
  /* fppowtf32.vhdl:5596:10  */
  always @(posedge clk)
    n1326 <= xsign_d5;
  /* fppowtf32.vhdl:5596:10  */
  always @(posedge clk)
    n1327 <= xsign_d6;
  /* fppowtf32.vhdl:5596:10  */
  always @(posedge clk)
    n1328 <= xexpfield;
  /* fppowtf32.vhdl:5596:10  */
  always @(posedge clk)
    n1329 <= e0;
  /* fppowtf32.vhdl:5596:10  */
  always @(posedge clk)
    n1330 <= e0_d1;
  /* fppowtf32.vhdl:5596:10  */
  always @(posedge clk)
    n1331 <= e0_d2;
  /* fppowtf32.vhdl:5596:10  */
  always @(posedge clk)
    n1332 <= e0_d3;
  /* fppowtf32.vhdl:5596:10  */
  always @(posedge clk)
    n1333 <= e0_d4;
  /* fppowtf32.vhdl:5596:10  */
  always @(posedge clk)
    n1334 <= e0_d5;
  /* fppowtf32.vhdl:5596:10  */
  always @(posedge clk)
    n1335 <= e0_d6;
  /* fppowtf32.vhdl:5596:10  */
  always @(posedge clk)
    n1336 <= e0_d7;
  /* fppowtf32.vhdl:5596:10  */
  always @(posedge clk)
    n1337 <= e0_d8;
  /* fppowtf32.vhdl:5596:10  */
  always @(posedge clk)
    n1338 <= e0_d9;
  /* fppowtf32.vhdl:5596:10  */
  always @(posedge clk)
    n1339 <= e0_d10;
  /* fppowtf32.vhdl:5596:10  */
  always @(posedge clk)
    n1340 <= e0_d11;
  /* fppowtf32.vhdl:5596:10  */
  always @(posedge clk)
    n1341 <= e0_d12;
  /* fppowtf32.vhdl:5596:10  */
  always @(posedge clk)
    n1342 <= e0_d13;
  /* fppowtf32.vhdl:5596:10  */
  always @(posedge clk)
    n1343 <= shiftval;
  /* fppowtf32.vhdl:5596:10  */
  always @(posedge clk)
    n1344 <= resultwillbeone;
  /* fppowtf32.vhdl:5596:10  */
  always @(posedge clk)
    n1345 <= maxshift;
  /* fppowtf32.vhdl:5596:10  */
  always @(posedge clk)
    n1346 <= maxshift_d1;
  /* fppowtf32.vhdl:5596:10  */
  always @(posedge clk)
    n1347 <= maxshift_d2;
  /* fppowtf32.vhdl:5596:10  */
  always @(posedge clk)
    n1348 <= maxshift_d3;
  /* fppowtf32.vhdl:5596:10  */
  always @(posedge clk)
    n1349 <= maxshift_d4;
  /* fppowtf32.vhdl:5596:10  */
  always @(posedge clk)
    n1350 <= maxshift_d5;
  /* fppowtf32.vhdl:5596:10  */
  always @(posedge clk)
    n1351 <= maxshift_d6;
  /* fppowtf32.vhdl:5596:10  */
  always @(posedge clk)
    n1352 <= maxshift_d7;
  /* fppowtf32.vhdl:5596:10  */
  always @(posedge clk)
    n1353 <= maxshift_d8;
  /* fppowtf32.vhdl:5596:10  */
  always @(posedge clk)
    n1354 <= maxshift_d9;
  /* fppowtf32.vhdl:5596:10  */
  always @(posedge clk)
    n1355 <= maxshift_d10;
  /* fppowtf32.vhdl:5596:10  */
  always @(posedge clk)
    n1356 <= maxshift_d11;
  /* fppowtf32.vhdl:5596:10  */
  always @(posedge clk)
    n1357 <= maxshift_d12;
  /* fppowtf32.vhdl:5596:10  */
  always @(posedge clk)
    n1358 <= maxshift_d13;
  /* fppowtf32.vhdl:5596:10  */
  always @(posedge clk)
    n1359 <= maxshift_d14;
  /* fppowtf32.vhdl:5596:10  */
  always @(posedge clk)
    n1360 <= k;
  /* fppowtf32.vhdl:5596:10  */
  always @(posedge clk)
    n1361 <= k_d1;
  /* fppowtf32.vhdl:5596:10  */
  always @(posedge clk)
    n1362 <= ofl1;
  /* fppowtf32.vhdl:5596:10  */
  always @(posedge clk)
    n1363 <= ofl1_d1;
  /* fppowtf32.vhdl:5596:10  */
  always @(posedge clk)
    n1364 <= ofl1_d2;
  /* fppowtf32.vhdl:5596:10  */
  always @(posedge clk)
    n1365 <= ofl1_d3;
  /* fppowtf32.vhdl:5596:10  */
  always @(posedge clk)
    n1366 <= ofl1_d4;
  /* fppowtf32.vhdl:5596:10  */
  always @(posedge clk)
    n1367 <= ofl3;
  /* fppowtf32.vhdl:5596:10  */
  always @(posedge clk)
    n1368 <= ofl3_d1;
  /* fppowtf32.vhdl:5596:10  */
  always @(posedge clk)
    n1369 <= ofl3_d2;
  /* fppowtf32.vhdl:5596:10  */
  always @(posedge clk)
    n1370 <= ofl3_d3;
  /* fppowtf32.vhdl:5596:10  */
  always @(posedge clk)
    n1371 <= ofl3_d4;
  /* fppowtf32.vhdl:5596:10  */
  always @(posedge clk)
    n1372 <= ofl3_d5;
  /* fppowtf32.vhdl:5596:10  */
  always @(posedge clk)
    n1373 <= ofl3_d6;
  /* fppowtf32.vhdl:5596:10  */
  always @(posedge clk)
    n1374 <= ufl2;
  /* fppowtf32.vhdl:5596:10  */
  always @(posedge clk)
    n1375 <= ufl2_d1;
  /* fppowtf32.vhdl:5596:10  */
  always @(posedge clk)
    n1376 <= ufl2_d2;
  /* fppowtf32.vhdl:5596:10  */
  always @(posedge clk)
    n1377 <= ufl2_d3;
  /* fppowtf32.vhdl:5596:10  */
  always @(posedge clk)
    n1378 <= ufl2_d4;
  /* fppowtf32.vhdl:5596:10  */
  always @(posedge clk)
    n1379 <= ufl2_d5;
  /* fppowtf32.vhdl:5596:10  */
  always @(posedge clk)
    n1380 <= ufl2_d6;
  /* fppowtf32.vhdl:5596:10  */
  always @(posedge clk)
    n1381 <= ufl3;
  /* fppowtf32.vhdl:5596:10  */
  always @(posedge clk)
    n1382 <= ufl3_d1;
  /* fppowtf32.vhdl:5596:10  */
  always @(posedge clk)
    n1383 <= ufl3_d2;
  /* fppowtf32.vhdl:5596:10  */
  always @(posedge clk)
    n1384 <= ufl3_d3;
  /* fppowtf32.vhdl:5596:10  */
  always @(posedge clk)
    n1385 <= ufl3_d4;
endmodule

module fpmult_8_20_uid62_freq500_uid63
  (input  clk,
   input  [30:0] x,
   input  [20:0] y,
   output [31:0] r);
  wire sign;
  wire sign_d1;
  wire sign_d2;
  wire [7:0] expx;
  wire [7:0] expx_d1;
  wire [7:0] expy;
  wire [7:0] expy_d1;
  wire [7:0] expy_d2;
  wire [7:0] expy_d3;
  wire [7:0] expy_d4;
  wire [7:0] expy_d5;
  wire [7:0] expy_d6;
  wire [7:0] expy_d7;
  wire [7:0] expy_d8;
  wire [7:0] expy_d9;
  wire [7:0] expy_d10;
  wire [7:0] expy_d11;
  wire [7:0] expy_d12;
  wire [9:0] expsumpresub;
  wire [9:0] expsumpresub_d1;
  wire [9:0] bias;
  wire [9:0] bias_d1;
  wire [9:0] bias_d2;
  wire [9:0] bias_d3;
  wire [9:0] bias_d4;
  wire [9:0] bias_d5;
  wire [9:0] bias_d6;
  wire [9:0] bias_d7;
  wire [9:0] bias_d8;
  wire [9:0] bias_d9;
  wire [9:0] bias_d10;
  wire [9:0] bias_d11;
  wire [9:0] bias_d12;
  wire [9:0] bias_d13;
  wire [9:0] expsum;
  wire [20:0] sigx;
  wire [10:0] sigy;
  wire [23:0] sigprod;
  wire [23:0] sigprod_d1;
  wire [3:0] excsel;
  wire [1:0] exc;
  wire [1:0] exc_d1;
  wire [1:0] exc_d2;
  wire norm;
  wire norm_d1;
  wire norm_d2;
  wire [9:0] exppostnorm;
  wire [23:0] sigprodext;
  wire [23:0] sigprodext_d1;
  wire [30:0] expsig;
  wire round;
  wire [30:0] expsigpostround;
  wire [1:0] excpostnorm;
  wire [1:0] finalexc;
  wire [20:0] y_d1;
  wire [20:0] y_d2;
  wire [20:0] y_d3;
  wire [20:0] y_d4;
  wire [20:0] y_d5;
  wire [20:0] y_d6;
  wire [20:0] y_d7;
  wire [20:0] y_d8;
  wire [20:0] y_d9;
  wire [20:0] y_d10;
  wire [20:0] y_d11;
  wire n981;
  wire n982;
  wire n983;
  wire [7:0] n984;
  wire [7:0] n985;
  wire [9:0] n987;
  wire [9:0] n989;
  wire [9:0] n990;
  wire [9:0] n992;
  wire [19:0] n993;
  wire [20:0] n995;
  wire [9:0] n996;
  wire [10:0] n998;
  wire [23:0] significandmultiplication_n999;
  wire [1:0] n1002;
  wire [1:0] n1003;
  wire [3:0] n1004;
  wire n1007;
  wire n1009;
  wire n1010;
  wire n1012;
  wire n1013;
  wire n1016;
  wire n1019;
  wire n1021;
  wire n1022;
  wire n1024;
  wire n1025;
  wire [2:0] n1027;
  reg [1:0] n1028;
  wire n1029;
  wire [9:0] n1031;
  wire [9:0] n1032;
  wire [22:0] n1033;
  wire [23:0] n1035;
  wire [23:0] n1036;
  wire [21:0] n1037;
  wire [23:0] n1039;
  wire [20:0] n1040;
  wire [30:0] n1041;
  localparam [30:0] n1043 = 31'b0000000000000000000000000000000;
  wire [30:0] roundingadder_n1044;
  wire [1:0] n1047;
  wire n1050;
  wire n1053;
  wire n1056;
  wire n1058;
  wire n1059;
  wire [2:0] n1061;
  reg [1:0] n1062;
  wire n1064;
  wire n1066;
  wire n1067;
  wire n1069;
  wire n1070;
  reg [1:0] n1071;
  wire [2:0] n1072;
  wire [28:0] n1073;
  wire [31:0] n1074;
  reg n1075;
  reg n1076;
  reg [7:0] n1077;
  reg [7:0] n1078;
  reg [7:0] n1079;
  reg [7:0] n1080;
  reg [7:0] n1081;
  reg [7:0] n1082;
  reg [7:0] n1083;
  reg [7:0] n1084;
  reg [7:0] n1085;
  reg [7:0] n1086;
  reg [7:0] n1087;
  reg [7:0] n1088;
  reg [7:0] n1089;
  reg [9:0] n1090;
  reg [9:0] n1091;
  reg [9:0] n1092;
  reg [9:0] n1093;
  reg [9:0] n1094;
  reg [9:0] n1095;
  reg [9:0] n1096;
  reg [9:0] n1097;
  reg [9:0] n1098;
  reg [9:0] n1099;
  reg [9:0] n1100;
  reg [9:0] n1101;
  reg [9:0] n1102;
  reg [9:0] n1103;
  reg [23:0] n1104;
  reg [1:0] n1105;
  reg [1:0] n1106;
  reg n1107;
  reg n1108;
  reg [23:0] n1109;
  reg [20:0] n1110;
  reg [20:0] n1111;
  reg [20:0] n1112;
  reg [20:0] n1113;
  reg [20:0] n1114;
  reg [20:0] n1115;
  reg [20:0] n1116;
  reg [20:0] n1117;
  reg [20:0] n1118;
  reg [20:0] n1119;
  reg [20:0] n1120;
  assign r = n1074; //(module output)
  /* fppowtf32.vhdl:4208:8  */
  assign sign = n983; // (signal)
  /* fppowtf32.vhdl:4208:14  */
  assign sign_d1 = n1075; // (signal)
  /* fppowtf32.vhdl:4208:23  */
  assign sign_d2 = n1076; // (signal)
  /* fppowtf32.vhdl:4210:8  */
  assign expx = n984; // (signal)
  /* fppowtf32.vhdl:4210:14  */
  assign expx_d1 = n1077; // (signal)
  /* fppowtf32.vhdl:4212:8  */
  assign expy = n985; // (signal)
  /* fppowtf32.vhdl:4212:14  */
  assign expy_d1 = n1078; // (signal)
  /* fppowtf32.vhdl:4212:23  */
  assign expy_d2 = n1079; // (signal)
  /* fppowtf32.vhdl:4212:32  */
  assign expy_d3 = n1080; // (signal)
  /* fppowtf32.vhdl:4212:41  */
  assign expy_d4 = n1081; // (signal)
  /* fppowtf32.vhdl:4212:50  */
  assign expy_d5 = n1082; // (signal)
  /* fppowtf32.vhdl:4212:59  */
  assign expy_d6 = n1083; // (signal)
  /* fppowtf32.vhdl:4212:68  */
  assign expy_d7 = n1084; // (signal)
  /* fppowtf32.vhdl:4212:77  */
  assign expy_d8 = n1085; // (signal)
  /* fppowtf32.vhdl:4212:86  */
  assign expy_d9 = n1086; // (signal)
  /* fppowtf32.vhdl:4212:95  */
  assign expy_d10 = n1087; // (signal)
  /* fppowtf32.vhdl:4212:105  */
  assign expy_d11 = n1088; // (signal)
  /* fppowtf32.vhdl:4212:115  */
  assign expy_d12 = n1089; // (signal)
  /* fppowtf32.vhdl:4214:8  */
  assign expsumpresub = n990; // (signal)
  /* fppowtf32.vhdl:4214:22  */
  assign expsumpresub_d1 = n1090; // (signal)
  /* fppowtf32.vhdl:4216:8  */
  assign bias = 10'b0001111111; // (signal)
  /* fppowtf32.vhdl:4216:14  */
  assign bias_d1 = n1091; // (signal)
  /* fppowtf32.vhdl:4216:23  */
  assign bias_d2 = n1092; // (signal)
  /* fppowtf32.vhdl:4216:32  */
  assign bias_d3 = n1093; // (signal)
  /* fppowtf32.vhdl:4216:41  */
  assign bias_d4 = n1094; // (signal)
  /* fppowtf32.vhdl:4216:50  */
  assign bias_d5 = n1095; // (signal)
  /* fppowtf32.vhdl:4216:59  */
  assign bias_d6 = n1096; // (signal)
  /* fppowtf32.vhdl:4216:68  */
  assign bias_d7 = n1097; // (signal)
  /* fppowtf32.vhdl:4216:77  */
  assign bias_d8 = n1098; // (signal)
  /* fppowtf32.vhdl:4216:86  */
  assign bias_d9 = n1099; // (signal)
  /* fppowtf32.vhdl:4216:95  */
  assign bias_d10 = n1100; // (signal)
  /* fppowtf32.vhdl:4216:105  */
  assign bias_d11 = n1101; // (signal)
  /* fppowtf32.vhdl:4216:115  */
  assign bias_d12 = n1102; // (signal)
  /* fppowtf32.vhdl:4216:125  */
  assign bias_d13 = n1103; // (signal)
  /* fppowtf32.vhdl:4218:8  */
  assign expsum = n992; // (signal)
  /* fppowtf32.vhdl:4220:8  */
  assign sigx = n995; // (signal)
  /* fppowtf32.vhdl:4222:8  */
  assign sigy = n998; // (signal)
  /* fppowtf32.vhdl:4224:8  */
  assign sigprod = significandmultiplication_n999; // (signal)
  /* fppowtf32.vhdl:4224:17  */
  assign sigprod_d1 = n1104; // (signal)
  /* fppowtf32.vhdl:4226:8  */
  assign excsel = n1004; // (signal)
  /* fppowtf32.vhdl:4228:8  */
  assign exc = n1028; // (signal)
  /* fppowtf32.vhdl:4228:13  */
  assign exc_d1 = n1105; // (signal)
  /* fppowtf32.vhdl:4228:21  */
  assign exc_d2 = n1106; // (signal)
  /* fppowtf32.vhdl:4230:8  */
  assign norm = n1029; // (signal)
  /* fppowtf32.vhdl:4230:14  */
  assign norm_d1 = n1107; // (signal)
  /* fppowtf32.vhdl:4230:23  */
  assign norm_d2 = n1108; // (signal)
  /* fppowtf32.vhdl:4232:8  */
  assign exppostnorm = n1032; // (signal)
  /* fppowtf32.vhdl:4234:8  */
  assign sigprodext = n1036; // (signal)
  /* fppowtf32.vhdl:4234:20  */
  assign sigprodext_d1 = n1109; // (signal)
  /* fppowtf32.vhdl:4236:8  */
  assign expsig = n1041; // (signal)
  /* fppowtf32.vhdl:4238:8  */
  assign round = 1'b1; // (signal)
  /* fppowtf32.vhdl:4240:8  */
  assign expsigpostround = roundingadder_n1044; // (signal)
  /* fppowtf32.vhdl:4242:8  */
  assign excpostnorm = n1062; // (signal)
  /* fppowtf32.vhdl:4244:8  */
  assign finalexc = n1071; // (signal)
  /* fppowtf32.vhdl:4246:8  */
  assign y_d1 = n1110; // (signal)
  /* fppowtf32.vhdl:4246:14  */
  assign y_d2 = n1111; // (signal)
  /* fppowtf32.vhdl:4246:20  */
  assign y_d3 = n1112; // (signal)
  /* fppowtf32.vhdl:4246:26  */
  assign y_d4 = n1113; // (signal)
  /* fppowtf32.vhdl:4246:32  */
  assign y_d5 = n1114; // (signal)
  /* fppowtf32.vhdl:4246:38  */
  assign y_d6 = n1115; // (signal)
  /* fppowtf32.vhdl:4246:44  */
  assign y_d7 = n1116; // (signal)
  /* fppowtf32.vhdl:4246:50  */
  assign y_d8 = n1117; // (signal)
  /* fppowtf32.vhdl:4246:56  */
  assign y_d9 = n1118; // (signal)
  /* fppowtf32.vhdl:4246:62  */
  assign y_d10 = n1119; // (signal)
  /* fppowtf32.vhdl:4246:69  */
  assign y_d11 = n1120; // (signal)
  /* fppowtf32.vhdl:4300:13  */
  assign n981 = x[28]; // extract
  /* fppowtf32.vhdl:4300:27  */
  assign n982 = y_d11[18]; // extract
  /* fppowtf32.vhdl:4300:18  */
  assign n983 = n981 ^ n982;
  /* fppowtf32.vhdl:4301:13  */
  assign n984 = x[27:20]; // extract
  /* fppowtf32.vhdl:4302:13  */
  assign n985 = y[17:10]; // extract
  /* fppowtf32.vhdl:4303:26  */
  assign n987 = {2'b00, expx_d1};
  /* fppowtf32.vhdl:4303:45  */
  assign n989 = {2'b00, expy_d12};
  /* fppowtf32.vhdl:4303:37  */
  assign n990 = n987 + n989;
  /* fppowtf32.vhdl:4305:30  */
  assign n992 = expsumpresub_d1 - bias_d13;
  /* fppowtf32.vhdl:4306:19  */
  assign n993 = x[19:0]; // extract
  /* fppowtf32.vhdl:4306:16  */
  assign n995 = {1'b1, n993};
  /* fppowtf32.vhdl:4307:19  */
  assign n996 = y[9:0]; // extract
  /* fppowtf32.vhdl:4307:16  */
  assign n998 = {1'b1, n996};
  /* fppowtf32.vhdl:4308:4  */
  intmultiplier_21x11_24_freq500_uid65 significandmultiplication (
    .clk(clk),
    .x(sigx),
    .y(sigy),
    .r(significandmultiplication_n999));
  /* fppowtf32.vhdl:4313:15  */
  assign n1002 = x[30:29]; // extract
  /* fppowtf32.vhdl:4313:37  */
  assign n1003 = y_d11[20:19]; // extract
  /* fppowtf32.vhdl:4313:30  */
  assign n1004 = {n1002, n1003};
  /* fppowtf32.vhdl:4315:16  */
  assign n1007 = excsel == 4'b0000;
  /* fppowtf32.vhdl:4315:29  */
  assign n1009 = excsel == 4'b0001;
  /* fppowtf32.vhdl:4315:29  */
  assign n1010 = n1007 | n1009;
  /* fppowtf32.vhdl:4315:38  */
  assign n1012 = excsel == 4'b0100;
  /* fppowtf32.vhdl:4315:38  */
  assign n1013 = n1010 | n1012;
  /* fppowtf32.vhdl:4316:16  */
  assign n1016 = excsel == 4'b0101;
  /* fppowtf32.vhdl:4317:16  */
  assign n1019 = excsel == 4'b0110;
  /* fppowtf32.vhdl:4317:28  */
  assign n1021 = excsel == 4'b1001;
  /* fppowtf32.vhdl:4317:28  */
  assign n1022 = n1019 | n1021;
  /* fppowtf32.vhdl:4317:37  */
  assign n1024 = excsel == 4'b1010;
  /* fppowtf32.vhdl:4317:37  */
  assign n1025 = n1022 | n1024;
  assign n1027 = {n1025, n1016, n1013};
  /* fppowtf32.vhdl:4314:4  */
  always @*
    case (n1027)
      3'b100: n1028 = 2'b10;
      3'b010: n1028 = 2'b01;
      3'b001: n1028 = 2'b00;
      default: n1028 = 2'b11;
    endcase
  /* fppowtf32.vhdl:4319:19  */
  assign n1029 = sigprod[23]; // extract
  /* fppowtf32.vhdl:4321:41  */
  assign n1031 = {9'b000000000, norm_d2};
  /* fppowtf32.vhdl:4321:26  */
  assign n1032 = expsum + n1031;
  /* fppowtf32.vhdl:4323:28  */
  assign n1033 = sigprod_d1[22:0]; // extract
  /* fppowtf32.vhdl:4323:42  */
  assign n1035 = {n1033, 1'b0};
  /* fppowtf32.vhdl:4323:48  */
  assign n1036 = norm_d1 ? n1035 : n1039;
  /* fppowtf32.vhdl:4324:36  */
  assign n1037 = sigprod_d1[21:0]; // extract
  /* fppowtf32.vhdl:4324:50  */
  assign n1039 = {n1037, 2'b00};
  /* fppowtf32.vhdl:4325:41  */
  assign n1040 = sigprodext_d1[23:3]; // extract
  /* fppowtf32.vhdl:4325:26  */
  assign n1041 = {exppostnorm, n1040};
  /* fppowtf32.vhdl:4327:4  */
  intadder_31_freq500_uid69 roundingadder (
    .clk(clk),
    .x(expsig),
    .y(n1043),
    .cin(round),
    .r(roundingadder_n1044));
  /* fppowtf32.vhdl:4333:24  */
  assign n1047 = expsigpostround[30:29]; // extract
  /* fppowtf32.vhdl:4334:26  */
  assign n1050 = n1047 == 2'b00;
  /* fppowtf32.vhdl:4335:49  */
  assign n1053 = n1047 == 2'b01;
  /* fppowtf32.vhdl:4336:49  */
  assign n1056 = n1047 == 2'b11;
  /* fppowtf32.vhdl:4336:58  */
  assign n1058 = n1047 == 2'b10;
  /* fppowtf32.vhdl:4336:58  */
  assign n1059 = n1056 | n1058;
  assign n1061 = {n1059, n1053, n1050};
  /* fppowtf32.vhdl:4333:4  */
  always @*
    case (n1061)
      3'b100: n1062 = 2'b00;
      3'b010: n1062 = 2'b10;
      3'b001: n1062 = 2'b01;
      default: n1062 = 2'b11;
    endcase
  /* fppowtf32.vhdl:4339:23  */
  assign n1064 = exc_d2 == 2'b11;
  /* fppowtf32.vhdl:4339:33  */
  assign n1066 = exc_d2 == 2'b10;
  /* fppowtf32.vhdl:4339:33  */
  assign n1067 = n1064 | n1066;
  /* fppowtf32.vhdl:4339:38  */
  assign n1069 = exc_d2 == 2'b00;
  /* fppowtf32.vhdl:4339:38  */
  assign n1070 = n1067 | n1069;
  /* fppowtf32.vhdl:4338:4  */
  always @*
    case (n1070)
      1'b1: n1071 = exc_d2;
      default: n1071 = excpostnorm;
    endcase
  /* fppowtf32.vhdl:4341:18  */
  assign n1072 = {finalexc, sign_d2};
  /* fppowtf32.vhdl:4341:45  */
  assign n1073 = expsigpostround[28:0]; // extract
  /* fppowtf32.vhdl:4341:28  */
  assign n1074 = {n1072, n1073};
  /* fppowtf32.vhdl:4251:10  */
  always @(posedge clk)
    n1075 <= sign;
  /* fppowtf32.vhdl:4251:10  */
  always @(posedge clk)
    n1076 <= sign_d1;
  /* fppowtf32.vhdl:4251:10  */
  always @(posedge clk)
    n1077 <= expx;
  /* fppowtf32.vhdl:4251:10  */
  always @(posedge clk)
    n1078 <= expy;
  /* fppowtf32.vhdl:4251:10  */
  always @(posedge clk)
    n1079 <= expy_d1;
  /* fppowtf32.vhdl:4251:10  */
  always @(posedge clk)
    n1080 <= expy_d2;
  /* fppowtf32.vhdl:4251:10  */
  always @(posedge clk)
    n1081 <= expy_d3;
  /* fppowtf32.vhdl:4251:10  */
  always @(posedge clk)
    n1082 <= expy_d4;
  /* fppowtf32.vhdl:4251:10  */
  always @(posedge clk)
    n1083 <= expy_d5;
  /* fppowtf32.vhdl:4251:10  */
  always @(posedge clk)
    n1084 <= expy_d6;
  /* fppowtf32.vhdl:4251:10  */
  always @(posedge clk)
    n1085 <= expy_d7;
  /* fppowtf32.vhdl:4251:10  */
  always @(posedge clk)
    n1086 <= expy_d8;
  /* fppowtf32.vhdl:4251:10  */
  always @(posedge clk)
    n1087 <= expy_d9;
  /* fppowtf32.vhdl:4251:10  */
  always @(posedge clk)
    n1088 <= expy_d10;
  /* fppowtf32.vhdl:4251:10  */
  always @(posedge clk)
    n1089 <= expy_d11;
  /* fppowtf32.vhdl:4251:10  */
  always @(posedge clk)
    n1090 <= expsumpresub;
  /* fppowtf32.vhdl:4251:10  */
  always @(posedge clk)
    n1091 <= bias;
  /* fppowtf32.vhdl:4251:10  */
  always @(posedge clk)
    n1092 <= bias_d1;
  /* fppowtf32.vhdl:4251:10  */
  always @(posedge clk)
    n1093 <= bias_d2;
  /* fppowtf32.vhdl:4251:10  */
  always @(posedge clk)
    n1094 <= bias_d3;
  /* fppowtf32.vhdl:4251:10  */
  always @(posedge clk)
    n1095 <= bias_d4;
  /* fppowtf32.vhdl:4251:10  */
  always @(posedge clk)
    n1096 <= bias_d5;
  /* fppowtf32.vhdl:4251:10  */
  always @(posedge clk)
    n1097 <= bias_d6;
  /* fppowtf32.vhdl:4251:10  */
  always @(posedge clk)
    n1098 <= bias_d7;
  /* fppowtf32.vhdl:4251:10  */
  always @(posedge clk)
    n1099 <= bias_d8;
  /* fppowtf32.vhdl:4251:10  */
  always @(posedge clk)
    n1100 <= bias_d9;
  /* fppowtf32.vhdl:4251:10  */
  always @(posedge clk)
    n1101 <= bias_d10;
  /* fppowtf32.vhdl:4251:10  */
  always @(posedge clk)
    n1102 <= bias_d11;
  /* fppowtf32.vhdl:4251:10  */
  always @(posedge clk)
    n1103 <= bias_d12;
  /* fppowtf32.vhdl:4251:10  */
  always @(posedge clk)
    n1104 <= sigprod;
  /* fppowtf32.vhdl:4251:10  */
  always @(posedge clk)
    n1105 <= exc;
  /* fppowtf32.vhdl:4251:10  */
  always @(posedge clk)
    n1106 <= exc_d1;
  /* fppowtf32.vhdl:4251:10  */
  always @(posedge clk)
    n1107 <= norm;
  /* fppowtf32.vhdl:4251:10  */
  always @(posedge clk)
    n1108 <= norm_d1;
  /* fppowtf32.vhdl:4251:10  */
  always @(posedge clk)
    n1109 <= sigprodext;
  /* fppowtf32.vhdl:4251:10  */
  always @(posedge clk)
    n1110 <= y;
  /* fppowtf32.vhdl:4251:10  */
  always @(posedge clk)
    n1111 <= y_d1;
  /* fppowtf32.vhdl:4251:10  */
  always @(posedge clk)
    n1112 <= y_d2;
  /* fppowtf32.vhdl:4251:10  */
  always @(posedge clk)
    n1113 <= y_d3;
  /* fppowtf32.vhdl:4251:10  */
  always @(posedge clk)
    n1114 <= y_d4;
  /* fppowtf32.vhdl:4251:10  */
  always @(posedge clk)
    n1115 <= y_d5;
  /* fppowtf32.vhdl:4251:10  */
  always @(posedge clk)
    n1116 <= y_d6;
  /* fppowtf32.vhdl:4251:10  */
  always @(posedge clk)
    n1117 <= y_d7;
  /* fppowtf32.vhdl:4251:10  */
  always @(posedge clk)
    n1118 <= y_d8;
  /* fppowtf32.vhdl:4251:10  */
  always @(posedge clk)
    n1119 <= y_d9;
  /* fppowtf32.vhdl:4251:10  */
  always @(posedge clk)
    n1120 <= y_d10;
endmodule

module fplogiterative_8_20_0_500_freq500_uid9
  (input  clk,
   input  [30:0] x,
   output [30:0] r);
  wire [2:0] xexnsgn;
  wire [2:0] xexnsgn_d1;
  wire [2:0] xexnsgn_d2;
  wire [2:0] xexnsgn_d3;
  wire [2:0] xexnsgn_d4;
  wire [2:0] xexnsgn_d5;
  wire [2:0] xexnsgn_d6;
  wire [2:0] xexnsgn_d7;
  wire [2:0] xexnsgn_d8;
  wire [2:0] xexnsgn_d9;
  wire [2:0] xexnsgn_d10;
  wire [2:0] xexnsgn_d11;
  wire firstbit;
  wire [21:0] y0;
  wire [21:0] y0_d1;
  wire [19:0] y0h;
  wire sr;
  wire sr_d1;
  wire sr_d2;
  wire sr_d3;
  wire sr_d4;
  wire sr_d5;
  wire sr_d6;
  wire sr_d7;
  wire sr_d8;
  wire sr_d9;
  wire sr_d10;
  wire sr_d11;
  wire [10:0] absz0;
  wire [7:0] e;
  wire [7:0] abse;
  wire eeqzero;
  wire eeqzero_d1;
  wire eeqzero_d2;
  wire eeqzero_d3;
  wire eeqzero_d4;
  wire [4:0] lzo;
  wire [4:0] lzo_d1;
  wire [4:0] lzo_d2;
  wire [4:0] lzo_d3;
  wire [4:0] pfinal_s;
  wire [4:0] pfinal_s_d1;
  wire [4:0] pfinal_s_d2;
  wire [4:0] pfinal_s_d3;
  wire [5:0] shiftval;
  wire [3:0] shiftvalinl;
  wire [3:0] shiftvalinr;
  wire dorr;
  wire dorr_d1;
  wire dorr_d2;
  wire \small ;
  wire small_d1;
  wire small_d2;
  wire small_d3;
  wire small_d4;
  wire small_d5;
  wire small_d6;
  wire small_d7;
  wire [21:0] small_absz0_normd_full;
  wire [10:0] small_absz0_normd;
  wire [10:0] small_absz0_normd_d1;
  wire [7:0] a0;
  wire [8:0] inva0;
  wire [8:0] inva0_d1;
  wire [8:0] inva0_copy16;
  wire [30:0] p0;
  wire [22:0] z1;
  wire [5:0] a1;
  wire [5:0] a1_d1;
  wire [16:0] b1;
  wire [22:0] zm1;
  wire [22:0] zm1_d1;
  wire [28:0] p1;
  wire [29:0] y1;
  wire [23:0] eiy1;
  wire [23:0] addxiter1;
  wire [23:0] eiypb1;
  wire [23:0] pp1;
  wire [23:0] z2;
  wire [23:0] zfinal;
  wire [23:0] zfinal_d1;
  wire [23:0] zfinal_d2;
  wire [14:0] squarerin;
  wire [29:0] z2o2_full;
  wire [29:0] z2o2_full_dummy;
  wire [11:0] z2o2_normal;
  wire [23:0] addfinallog1py;
  wire [23:0] log1p_normal;
  wire [34:0] l0;
  wire [34:0] l0_copy28;
  wire [34:0] s1;
  wire [28:0] l1;
  wire [28:0] l1_copy31;
  wire [34:0] sopx1;
  wire [34:0] s2;
  wire [34:0] almostlog;
  wire [34:0] adderlogf_normaly;
  wire [34:0] logf_normal;
  wire [31:0] abselog2;
  wire [42:0] abselog2_pad;
  wire [42:0] logf_normal_pad;
  wire [42:0] lnaddx;
  wire [42:0] lnaddy;
  wire [42:0] log_normal;
  wire [34:0] log_normal_normd;
  wire [4:0] e_normal;
  wire [14:0] z2o2_small_bs;
  wire [28:0] z2o2_small_s;
  wire [25:0] z2o2_small;
  wire [25:0] z_small;
  wire [25:0] log_smally;
  wire nsrcin;
  wire [25:0] log_small;
  wire [1:0] e0_sub;
  wire ufl;
  wire ufl_d1;
  wire ufl_d2;
  wire ufl_d3;
  wire ufl_d4;
  wire ufl_d5;
  wire ufl_d6;
  wire ufl_d7;
  wire ufl_d8;
  wire ufl_d9;
  wire ufl_d10;
  wire ufl_d11;
  wire [7:0] e_small;
  wire [7:0] e_small_d1;
  wire [7:0] e_small_d2;
  wire [7:0] e_small_d3;
  wire [7:0] e_small_d4;
  wire [23:0] log_small_normd;
  wire [23:0] log_small_normd_d1;
  wire [23:0] log_small_normd_d2;
  wire [23:0] log_small_normd_d3;
  wire [23:0] log_small_normd_d4;
  wire [23:0] log_small_normd_d5;
  wire [7:0] e0offset;
  wire [7:0] e0offset_d1;
  wire [7:0] e0offset_d2;
  wire [7:0] e0offset_d3;
  wire [7:0] e0offset_d4;
  wire [7:0] e0offset_d5;
  wire [7:0] e0offset_d6;
  wire [7:0] e0offset_d7;
  wire [7:0] e0offset_d8;
  wire [7:0] e0offset_d9;
  wire [7:0] e0offset_d10;
  wire [7:0] er;
  wire [7:0] er_d1;
  wire [23:0] log_g;
  wire round;
  wire [27:0] frax;
  wire [27:0] fray;
  wire [27:0] efr;
  wire [2:0] rexn;
  wire [2:0] n602;
  wire n603;
  wire [19:0] n604;
  wire [20:0] n606;
  wire [21:0] n608;
  wire n609;
  wire [21:0] n610;
  wire [19:0] n611;
  wire [21:0] n613;
  wire [19:0] n614;
  wire [7:0] n616;
  wire n618;
  wire n619;
  wire n620;
  wire n621;
  wire [10:0] n622;
  wire n623;
  wire [10:0] n624;
  wire [10:0] n625;
  wire [10:0] n627;
  wire [7:0] n628;
  wire n629;
  wire [7:0] n631;
  wire [7:0] n632;
  wire [7:0] n634;
  wire [7:0] n635;
  wire n638;
  wire n639;
  wire [4:0] lzoc1_n641;
  wire [5:0] n646;
  wire [5:0] n648;
  wire [5:0] n649;
  wire [3:0] n650;
  wire [3:0] n651;
  wire n652;
  wire n653;
  wire n654;
  wire [21:0] small_lshift_n655;
  wire [10:0] n658;
  wire [7:0] n659;
  wire [8:0] inva0table_n660;
  wire [30:0] n663;
  wire [30:0] n664;
  wire [30:0] n665;
  wire [22:0] n666;
  wire [5:0] n667;
  wire [16:0] n668;
  wire [28:0] n669;
  wire [28:0] n670;
  wire [28:0] n671;
  wire [29:0] n673;
  wire [23:0] n674;
  wire n675;
  wire [23:0] n676;
  wire [22:0] n677;
  wire [23:0] n679;
  wire [17:0] n681;
  wire [23:0] n683;
  localparam n684 = 1'b0;
  wire [23:0] additer1_1_n685;
  wire [22:0] n688;
  wire [22:0] n689;
  wire [23:0] n691;
  localparam n692 = 1'b1;
  wire [23:0] additer2_1_n693;
  wire [14:0] n696;
  wire [14:0] n697;
  wire [14:0] n699;
  wire [29:0] n700;
  wire [29:0] n701;
  wire [29:0] n702;
  wire [11:0] n703;
  wire [11:0] n704;
  wire [23:0] n706;
  localparam n707 = 1'b1;
  wire [23:0] addfinallog1p_normaladder_n708;
  wire [34:0] logtable0_n711;
  wire [28:0] logtable1_n714;
  wire [34:0] n718;
  localparam n719 = 1'b0;
  wire [34:0] adders1_n720;
  wire [34:0] n724;
  localparam n725 = 1'b0;
  wire [34:0] adderlogf_normal_n726;
  wire [31:0] mullog2_n729;
  wire [42:0] n733;
  wire n734;
  wire n735;
  wire n736;
  wire n737;
  wire n738;
  wire n739;
  wire n740;
  wire n741;
  wire [3:0] n742;
  wire [3:0] n743;
  wire [7:0] n744;
  wire [42:0] n745;
  wire n746;
  wire [42:0] n747;
  wire [42:0] n748;
  wire [42:0] lnadder_n749;
  wire [4:0] final_norm_n752;
  wire [34:0] final_norm_n753;
  wire [14:0] n758;
  wire [28:0] ao_rshift_n759;
  wire [14:0] n762;
  wire [25:0] n764;
  wire [25:0] n766;
  wire [25:0] n767;
  wire [25:0] n768;
  wire n769;
  wire [25:0] log_small_adder_n770;
  wire n774;
  wire [1:0] n775;
  wire [1:0] n777;
  wire n779;
  wire [1:0] n780;
  wire [7:0] n784;
  wire [7:0] n786;
  wire [7:0] n787;
  wire [23:0] n788;
  wire n789;
  wire [23:0] n790;
  wire [23:0] n791;
  wire n792;
  wire [23:0] n793;
  wire [23:0] n794;
  wire [7:0] n796;
  wire [7:0] n798;
  wire [7:0] n799;
  wire [22:0] n800;
  wire [23:0] n802;
  wire [23:0] n803;
  wire [23:0] n804;
  wire n805;
  wire [19:0] n806;
  wire [27:0] n807;
  wire [27:0] n809;
  localparam n810 = 1'b0;
  wire [27:0] finalroundadder_n811;
  wire n815;
  wire n816;
  wire n817;
  wire n818;
  wire n819;
  wire n820;
  wire n821;
  wire n822;
  wire n823;
  wire [2:0] n824;
  wire [1:0] n826;
  wire n828;
  wire [2:0] n829;
  wire [1:0] n831;
  wire n833;
  wire [2:0] n834;
  wire [2:0] n836;
  wire n837;
  wire n838;
  wire n839;
  wire n840;
  wire n841;
  wire n842;
  wire n843;
  wire n844;
  wire n845;
  wire n846;
  wire [2:0] n847;
  wire [2:0] n849;
  wire [30:0] n850;
  reg [2:0] n851;
  reg [2:0] n852;
  reg [2:0] n853;
  reg [2:0] n854;
  reg [2:0] n855;
  reg [2:0] n856;
  reg [2:0] n857;
  reg [2:0] n858;
  reg [2:0] n859;
  reg [2:0] n860;
  reg [2:0] n861;
  reg [21:0] n862;
  reg n863;
  reg n864;
  reg n865;
  reg n866;
  reg n867;
  reg n868;
  reg n869;
  reg n870;
  reg n871;
  reg n872;
  reg n873;
  reg n874;
  reg n875;
  reg n876;
  reg n877;
  reg [4:0] n878;
  reg [4:0] n879;
  reg [4:0] n880;
  reg [4:0] n881;
  reg [4:0] n882;
  reg [4:0] n883;
  reg n884;
  reg n885;
  reg n886;
  reg n887;
  reg n888;
  reg n889;
  reg n890;
  reg n891;
  reg n892;
  reg [10:0] n893;
  reg [8:0] n894;
  reg [5:0] n895;
  reg [22:0] n896;
  reg [23:0] n897;
  reg [23:0] n898;
  reg n899;
  reg n900;
  reg n901;
  reg n902;
  reg n903;
  reg n904;
  reg n905;
  reg n906;
  reg n907;
  reg n908;
  reg n909;
  reg [7:0] n910;
  reg [7:0] n911;
  reg [7:0] n912;
  reg [7:0] n913;
  reg [23:0] n914;
  reg [23:0] n915;
  reg [23:0] n916;
  reg [23:0] n917;
  reg [23:0] n918;
  reg [7:0] n919;
  reg [7:0] n920;
  reg [7:0] n921;
  reg [7:0] n922;
  reg [7:0] n923;
  reg [7:0] n924;
  reg [7:0] n925;
  reg [7:0] n926;
  reg [7:0] n927;
  reg [7:0] n928;
  reg [7:0] n929;
  assign r = n850; //(module output)
  /* fppowtf32.vhdl:3604:8  */
  assign xexnsgn = n602; // (signal)
  /* fppowtf32.vhdl:3604:17  */
  assign xexnsgn_d1 = n851; // (signal)
  /* fppowtf32.vhdl:3604:29  */
  assign xexnsgn_d2 = n852; // (signal)
  /* fppowtf32.vhdl:3604:41  */
  assign xexnsgn_d3 = n853; // (signal)
  /* fppowtf32.vhdl:3604:53  */
  assign xexnsgn_d4 = n854; // (signal)
  /* fppowtf32.vhdl:3604:65  */
  assign xexnsgn_d5 = n855; // (signal)
  /* fppowtf32.vhdl:3604:77  */
  assign xexnsgn_d6 = n856; // (signal)
  /* fppowtf32.vhdl:3604:89  */
  assign xexnsgn_d7 = n857; // (signal)
  /* fppowtf32.vhdl:3604:101  */
  assign xexnsgn_d8 = n858; // (signal)
  /* fppowtf32.vhdl:3604:113  */
  assign xexnsgn_d9 = n859; // (signal)
  /* fppowtf32.vhdl:3604:125  */
  assign xexnsgn_d10 = n860; // (signal)
  /* fppowtf32.vhdl:3604:138  */
  assign xexnsgn_d11 = n861; // (signal)
  /* fppowtf32.vhdl:3606:8  */
  assign firstbit = n603; // (signal)
  /* fppowtf32.vhdl:3608:8  */
  assign y0 = n610; // (signal)
  /* fppowtf32.vhdl:3608:12  */
  assign y0_d1 = n862; // (signal)
  /* fppowtf32.vhdl:3610:8  */
  assign y0h = n614; // (signal)
  /* fppowtf32.vhdl:3612:8  */
  assign sr = n619; // (signal)
  /* fppowtf32.vhdl:3612:12  */
  assign sr_d1 = n863; // (signal)
  /* fppowtf32.vhdl:3612:19  */
  assign sr_d2 = n864; // (signal)
  /* fppowtf32.vhdl:3612:26  */
  assign sr_d3 = n865; // (signal)
  /* fppowtf32.vhdl:3612:33  */
  assign sr_d4 = n866; // (signal)
  /* fppowtf32.vhdl:3612:40  */
  assign sr_d5 = n867; // (signal)
  /* fppowtf32.vhdl:3612:47  */
  assign sr_d6 = n868; // (signal)
  /* fppowtf32.vhdl:3612:54  */
  assign sr_d7 = n869; // (signal)
  /* fppowtf32.vhdl:3612:61  */
  assign sr_d8 = n870; // (signal)
  /* fppowtf32.vhdl:3612:68  */
  assign sr_d9 = n871; // (signal)
  /* fppowtf32.vhdl:3612:75  */
  assign sr_d10 = n872; // (signal)
  /* fppowtf32.vhdl:3612:83  */
  assign sr_d11 = n873; // (signal)
  /* fppowtf32.vhdl:3614:8  */
  assign absz0 = n624; // (signal)
  /* fppowtf32.vhdl:3616:8  */
  assign e = n632; // (signal)
  /* fppowtf32.vhdl:3618:8  */
  assign abse = n635; // (signal)
  /* fppowtf32.vhdl:3620:8  */
  assign eeqzero = n639; // (signal)
  /* fppowtf32.vhdl:3620:17  */
  assign eeqzero_d1 = n874; // (signal)
  /* fppowtf32.vhdl:3620:29  */
  assign eeqzero_d2 = n875; // (signal)
  /* fppowtf32.vhdl:3620:41  */
  assign eeqzero_d3 = n876; // (signal)
  /* fppowtf32.vhdl:3620:53  */
  assign eeqzero_d4 = n877; // (signal)
  /* fppowtf32.vhdl:3622:8  */
  assign lzo = lzoc1_n641; // (signal)
  /* fppowtf32.vhdl:3622:13  */
  assign lzo_d1 = n878; // (signal)
  /* fppowtf32.vhdl:3622:21  */
  assign lzo_d2 = n879; // (signal)
  /* fppowtf32.vhdl:3622:29  */
  assign lzo_d3 = n880; // (signal)
  /* fppowtf32.vhdl:3624:8  */
  assign pfinal_s = 5'b01011; // (signal)
  /* fppowtf32.vhdl:3624:18  */
  assign pfinal_s_d1 = n881; // (signal)
  /* fppowtf32.vhdl:3624:31  */
  assign pfinal_s_d2 = n882; // (signal)
  /* fppowtf32.vhdl:3624:44  */
  assign pfinal_s_d3 = n883; // (signal)
  /* fppowtf32.vhdl:3626:8  */
  assign shiftval = n649; // (signal)
  /* fppowtf32.vhdl:3628:8  */
  assign shiftvalinl = n650; // (signal)
  /* fppowtf32.vhdl:3630:8  */
  assign shiftvalinr = n651; // (signal)
  /* fppowtf32.vhdl:3632:8  */
  assign dorr = n652; // (signal)
  /* fppowtf32.vhdl:3632:14  */
  assign dorr_d1 = n884; // (signal)
  /* fppowtf32.vhdl:3632:23  */
  assign dorr_d2 = n885; // (signal)
  /* fppowtf32.vhdl:3634:8  */
  assign \small  = n654; // (signal)
  /* fppowtf32.vhdl:3634:15  */
  assign small_d1 = n886; // (signal)
  /* fppowtf32.vhdl:3634:25  */
  assign small_d2 = n887; // (signal)
  /* fppowtf32.vhdl:3634:35  */
  assign small_d3 = n888; // (signal)
  /* fppowtf32.vhdl:3634:45  */
  assign small_d4 = n889; // (signal)
  /* fppowtf32.vhdl:3634:55  */
  assign small_d5 = n890; // (signal)
  /* fppowtf32.vhdl:3634:65  */
  assign small_d6 = n891; // (signal)
  /* fppowtf32.vhdl:3634:75  */
  assign small_d7 = n892; // (signal)
  /* fppowtf32.vhdl:3636:8  */
  assign small_absz0_normd_full = small_lshift_n655; // (signal)
  /* fppowtf32.vhdl:3638:8  */
  assign small_absz0_normd = n658; // (signal)
  /* fppowtf32.vhdl:3638:27  */
  assign small_absz0_normd_d1 = n893; // (signal)
  /* fppowtf32.vhdl:3640:8  */
  assign a0 = n659; // (signal)
  /* fppowtf32.vhdl:3642:8  */
  assign inva0 = inva0_copy16; // (signal)
  /* fppowtf32.vhdl:3642:15  */
  assign inva0_d1 = n894; // (signal)
  /* fppowtf32.vhdl:3644:8  */
  assign inva0_copy16 = inva0table_n660; // (signal)
  /* fppowtf32.vhdl:3646:8  */
  assign p0 = n665; // (signal)
  /* fppowtf32.vhdl:3648:8  */
  assign z1 = n666; // (signal)
  /* fppowtf32.vhdl:3650:8  */
  assign a1 = n667; // (signal)
  /* fppowtf32.vhdl:3650:12  */
  assign a1_d1 = n895; // (signal)
  /* fppowtf32.vhdl:3652:8  */
  assign b1 = n668; // (signal)
  /* fppowtf32.vhdl:3654:8  */
  assign zm1 = z1; // (signal)
  /* fppowtf32.vhdl:3654:13  */
  assign zm1_d1 = n896; // (signal)
  /* fppowtf32.vhdl:3656:8  */
  assign p1 = n671; // (signal)
  /* fppowtf32.vhdl:3658:8  */
  assign y1 = n673; // (signal)
  /* fppowtf32.vhdl:3660:8  */
  assign eiy1 = n676; // (signal)
  /* fppowtf32.vhdl:3662:8  */
  assign addxiter1 = n683; // (signal)
  /* fppowtf32.vhdl:3664:8  */
  assign eiypb1 = additer1_1_n685; // (signal)
  /* fppowtf32.vhdl:3666:8  */
  assign pp1 = n691; // (signal)
  /* fppowtf32.vhdl:3668:8  */
  assign z2 = additer2_1_n693; // (signal)
  /* fppowtf32.vhdl:3670:8  */
  assign zfinal = z2; // (signal)
  /* fppowtf32.vhdl:3670:16  */
  assign zfinal_d1 = n897; // (signal)
  /* fppowtf32.vhdl:3670:27  */
  assign zfinal_d2 = n898; // (signal)
  /* fppowtf32.vhdl:3672:8  */
  assign squarerin = n697; // (signal)
  /* fppowtf32.vhdl:3674:8  */
  assign z2o2_full = n702; // (signal)
  /* fppowtf32.vhdl:3676:8  */
  assign z2o2_full_dummy = z2o2_full; // (signal)
  /* fppowtf32.vhdl:3678:8  */
  assign z2o2_normal = n703; // (signal)
  /* fppowtf32.vhdl:3680:8  */
  assign addfinallog1py = n706; // (signal)
  /* fppowtf32.vhdl:3682:8  */
  assign log1p_normal = addfinallog1p_normaladder_n708; // (signal)
  /* fppowtf32.vhdl:3684:8  */
  assign l0 = l0_copy28; // (signal)
  /* fppowtf32.vhdl:3686:8  */
  assign l0_copy28 = logtable0_n711; // (signal)
  /* fppowtf32.vhdl:3688:8  */
  assign s1 = l0; // (signal)
  /* fppowtf32.vhdl:3690:8  */
  assign l1 = l1_copy31; // (signal)
  /* fppowtf32.vhdl:3692:8  */
  assign l1_copy31 = logtable1_n714; // (signal)
  /* fppowtf32.vhdl:3694:8  */
  assign sopx1 = n718; // (signal)
  /* fppowtf32.vhdl:3696:8  */
  assign s2 = adders1_n720; // (signal)
  /* fppowtf32.vhdl:3698:8  */
  assign almostlog = s2; // (signal)
  /* fppowtf32.vhdl:3700:8  */
  assign adderlogf_normaly = n724; // (signal)
  /* fppowtf32.vhdl:3702:8  */
  assign logf_normal = adderlogf_normal_n726; // (signal)
  /* fppowtf32.vhdl:3704:8  */
  assign abselog2 = mullog2_n729; // (signal)
  /* fppowtf32.vhdl:3706:8  */
  assign abselog2_pad = n733; // (signal)
  /* fppowtf32.vhdl:3708:8  */
  assign logf_normal_pad = n745; // (signal)
  /* fppowtf32.vhdl:3710:8  */
  assign lnaddx = abselog2_pad; // (signal)
  /* fppowtf32.vhdl:3712:8  */
  assign lnaddy = n747; // (signal)
  /* fppowtf32.vhdl:3714:8  */
  assign log_normal = lnadder_n749; // (signal)
  /* fppowtf32.vhdl:3716:8  */
  assign log_normal_normd = final_norm_n753; // (signal)
  /* fppowtf32.vhdl:3718:8  */
  assign e_normal = final_norm_n752; // (signal)
  /* fppowtf32.vhdl:3720:8  */
  assign z2o2_small_bs = n758; // (signal)
  /* fppowtf32.vhdl:3722:8  */
  assign z2o2_small_s = ao_rshift_n759; // (signal)
  /* fppowtf32.vhdl:3724:8  */
  assign z2o2_small = n764; // (signal)
  /* fppowtf32.vhdl:3726:8  */
  assign z_small = n766; // (signal)
  /* fppowtf32.vhdl:3728:8  */
  assign log_smally = n767; // (signal)
  /* fppowtf32.vhdl:3730:8  */
  assign nsrcin = n769; // (signal)
  /* fppowtf32.vhdl:3732:8  */
  assign log_small = log_small_adder_n770; // (signal)
  /* fppowtf32.vhdl:3734:8  */
  assign e0_sub = n775; // (signal)
  /* fppowtf32.vhdl:3736:8  */
  assign ufl = 1'b0; // (signal)
  /* fppowtf32.vhdl:3736:13  */
  assign ufl_d1 = n899; // (signal)
  /* fppowtf32.vhdl:3736:21  */
  assign ufl_d2 = n900; // (signal)
  /* fppowtf32.vhdl:3736:29  */
  assign ufl_d3 = n901; // (signal)
  /* fppowtf32.vhdl:3736:37  */
  assign ufl_d4 = n902; // (signal)
  /* fppowtf32.vhdl:3736:45  */
  assign ufl_d5 = n903; // (signal)
  /* fppowtf32.vhdl:3736:53  */
  assign ufl_d6 = n904; // (signal)
  /* fppowtf32.vhdl:3736:61  */
  assign ufl_d7 = n905; // (signal)
  /* fppowtf32.vhdl:3736:69  */
  assign ufl_d8 = n906; // (signal)
  /* fppowtf32.vhdl:3736:77  */
  assign ufl_d9 = n907; // (signal)
  /* fppowtf32.vhdl:3736:85  */
  assign ufl_d10 = n908; // (signal)
  /* fppowtf32.vhdl:3736:94  */
  assign ufl_d11 = n909; // (signal)
  /* fppowtf32.vhdl:3738:8  */
  assign e_small = n787; // (signal)
  /* fppowtf32.vhdl:3738:17  */
  assign e_small_d1 = n910; // (signal)
  /* fppowtf32.vhdl:3738:29  */
  assign e_small_d2 = n911; // (signal)
  /* fppowtf32.vhdl:3738:41  */
  assign e_small_d3 = n912; // (signal)
  /* fppowtf32.vhdl:3738:53  */
  assign e_small_d4 = n913; // (signal)
  /* fppowtf32.vhdl:3740:8  */
  assign log_small_normd = n790; // (signal)
  /* fppowtf32.vhdl:3740:25  */
  assign log_small_normd_d1 = n914; // (signal)
  /* fppowtf32.vhdl:3740:45  */
  assign log_small_normd_d2 = n915; // (signal)
  /* fppowtf32.vhdl:3740:65  */
  assign log_small_normd_d3 = n916; // (signal)
  /* fppowtf32.vhdl:3740:85  */
  assign log_small_normd_d4 = n917; // (signal)
  /* fppowtf32.vhdl:3740:105  */
  assign log_small_normd_d5 = n918; // (signal)
  /* fppowtf32.vhdl:3742:8  */
  assign e0offset = 8'b10000110; // (signal)
  /* fppowtf32.vhdl:3742:18  */
  assign e0offset_d1 = n919; // (signal)
  /* fppowtf32.vhdl:3742:31  */
  assign e0offset_d2 = n920; // (signal)
  /* fppowtf32.vhdl:3742:44  */
  assign e0offset_d3 = n921; // (signal)
  /* fppowtf32.vhdl:3742:57  */
  assign e0offset_d4 = n922; // (signal)
  /* fppowtf32.vhdl:3742:70  */
  assign e0offset_d5 = n923; // (signal)
  /* fppowtf32.vhdl:3742:83  */
  assign e0offset_d6 = n924; // (signal)
  /* fppowtf32.vhdl:3742:96  */
  assign e0offset_d7 = n925; // (signal)
  /* fppowtf32.vhdl:3742:109  */
  assign e0offset_d8 = n926; // (signal)
  /* fppowtf32.vhdl:3742:122  */
  assign e0offset_d9 = n927; // (signal)
  /* fppowtf32.vhdl:3742:135  */
  assign e0offset_d10 = n928; // (signal)
  /* fppowtf32.vhdl:3744:8  */
  assign er = n796; // (signal)
  /* fppowtf32.vhdl:3744:12  */
  assign er_d1 = n929; // (signal)
  /* fppowtf32.vhdl:3746:8  */
  assign log_g = n803; // (signal)
  /* fppowtf32.vhdl:3748:8  */
  assign round = n805; // (signal)
  /* fppowtf32.vhdl:3750:8  */
  assign frax = n807; // (signal)
  /* fppowtf32.vhdl:3752:8  */
  assign fray = n809; // (signal)
  /* fppowtf32.vhdl:3754:8  */
  assign efr = finalroundadder_n811; // (signal)
  /* fppowtf32.vhdl:3756:8  */
  assign rexn = n824; // (signal)
  /* fppowtf32.vhdl:3850:17  */
  assign n602 = x[30:28]; // extract
  /* fppowtf32.vhdl:3851:18  */
  assign n603 = x[19]; // extract
  /* fppowtf32.vhdl:3852:17  */
  assign n604 = x[19:0]; // extract
  /* fppowtf32.vhdl:3852:14  */
  assign n606 = {1'b1, n604};
  /* fppowtf32.vhdl:3852:33  */
  assign n608 = {n606, 1'b0};
  /* fppowtf32.vhdl:3852:53  */
  assign n609 = ~firstbit;
  /* fppowtf32.vhdl:3852:39  */
  assign n610 = n609 ? n608 : n613;
  /* fppowtf32.vhdl:3852:72  */
  assign n611 = x[19:0]; // extract
  /* fppowtf32.vhdl:3852:69  */
  assign n613 = {2'b01, n611};
  /* fppowtf32.vhdl:3853:13  */
  assign n614 = y0[20:1]; // extract
  /* fppowtf32.vhdl:3855:24  */
  assign n616 = x[27:20]; // extract
  /* fppowtf32.vhdl:3855:44  */
  assign n618 = n616 == 8'b01111111;
  /* fppowtf32.vhdl:3855:16  */
  assign n619 = n618 ? 1'b0 : n621;
  /* fppowtf32.vhdl:3856:16  */
  assign n620 = x[27]; // extract
  /* fppowtf32.vhdl:3856:11  */
  assign n621 = ~n620;
  /* fppowtf32.vhdl:3857:17  */
  assign n622 = y0[10:0]; // extract
  /* fppowtf32.vhdl:3857:57  */
  assign n623 = ~sr;
  /* fppowtf32.vhdl:3857:49  */
  assign n624 = n623 ? n622 : n627;
  /* fppowtf32.vhdl:3858:49  */
  assign n625 = y0[10:0]; // extract
  /* fppowtf32.vhdl:3858:45  */
  assign n627 = 11'b00000000000 - n625;
  /* fppowtf32.vhdl:3859:11  */
  assign n628 = x[27:20]; // extract
  /* fppowtf32.vhdl:3859:67  */
  assign n629 = ~firstbit;
  /* fppowtf32.vhdl:3859:64  */
  assign n631 = {7'b0111111, n629};
  /* fppowtf32.vhdl:3859:32  */
  assign n632 = n628 - n631;
  /* fppowtf32.vhdl:3860:36  */
  assign n634 = 8'b00000000 - e;
  /* fppowtf32.vhdl:3860:43  */
  assign n635 = sr ? n634 : e;
  /* fppowtf32.vhdl:3861:25  */
  assign n638 = e == 8'b00000000;
  /* fppowtf32.vhdl:3861:19  */
  assign n639 = n638 ? 1'b1 : 1'b0;
  /* fppowtf32.vhdl:3862:4  */
  lzoc_20_freq500_uid11 lzoc1 (
    .clk(clk),
    .i(y0h),
    .ozb(firstbit),
    .o(lzoc1_n641));
  /* fppowtf32.vhdl:3868:21  */
  assign n646 = {1'b0, lzo};
  /* fppowtf32.vhdl:3868:35  */
  assign n648 = {1'b0, pfinal_s_d3};
  /* fppowtf32.vhdl:3868:28  */
  assign n649 = n646 - n648;
  /* fppowtf32.vhdl:3869:27  */
  assign n650 = shiftval[3:0]; // extract
  /* fppowtf32.vhdl:3870:27  */
  assign n651 = shiftval[3:0]; // extract
  /* fppowtf32.vhdl:3871:20  */
  assign n652 = shiftval[5]; // extract
  /* fppowtf32.vhdl:3872:28  */
  assign n653 = ~dorr_d1;
  /* fppowtf32.vhdl:3872:24  */
  assign n654 = eeqzero_d4 & n653;
  /* fppowtf32.vhdl:3874:4  */
  leftshifter11_by_max_11_freq500_uid13 small_lshift (
    .clk(clk),
    .x(absz0),
    .s(shiftvalinl),
    .r(small_lshift_n655));
  /* fppowtf32.vhdl:3879:47  */
  assign n658 = small_absz0_normd_full[10:0]; // extract
  /* fppowtf32.vhdl:3881:11  */
  assign n659 = x[19:12]; // extract
  /* fppowtf32.vhdl:3883:4  */
  inva0table_freq500_uid15 inva0table (
    .x(a0),
    .y(inva0table_n660));
  /* fppowtf32.vhdl:3887:19  */
  assign n663 = {22'b0, inva0_d1};  //  uext
  /* fppowtf32.vhdl:3887:19  */
  assign n664 = {9'b0, y0_d1};  //  uext
  /* fppowtf32.vhdl:3887:19  */
  assign n665 = n663 * n664; // umul
  /* fppowtf32.vhdl:3889:12  */
  assign n666 = p0[22:0]; // extract
  /* fppowtf32.vhdl:3891:12  */
  assign n667 = z1[22:17]; // extract
  /* fppowtf32.vhdl:3892:12  */
  assign n668 = z1[16:0]; // extract
  /* fppowtf32.vhdl:3894:15  */
  assign n669 = {23'b0, a1_d1};  //  uext
  /* fppowtf32.vhdl:3894:15  */
  assign n670 = {6'b0, zm1_d1};  //  uext
  /* fppowtf32.vhdl:3894:15  */
  assign n671 = n669 * n670; // umul
  /* fppowtf32.vhdl:3895:36  */
  assign n673 = {7'b1000000, z1};
  /* fppowtf32.vhdl:3896:14  */
  assign n674 = y1[29:6]; // extract
  /* fppowtf32.vhdl:3896:36  */
  assign n675 = a1[5]; // extract
  /* fppowtf32.vhdl:3896:29  */
  assign n676 = n675 ? n674 : n679;
  /* fppowtf32.vhdl:3897:20  */
  assign n677 = y1[29:7]; // extract
  /* fppowtf32.vhdl:3897:16  */
  assign n679 = {1'b0, n677};
  /* fppowtf32.vhdl:3898:21  */
  assign n681 = {1'b0, b1};
  /* fppowtf32.vhdl:3898:26  */
  assign n683 = {n681, 6'b000000};
  /* fppowtf32.vhdl:3899:4  */
  intadder_24_freq500_uid19 additer1_1 (
    .clk(clk),
    .x(addxiter1),
    .y(eiy1),
    .cin(n684),
    .r(additer1_1_n685));
  /* fppowtf32.vhdl:3905:39  */
  assign n688 = p1[28:6]; // extract
  /* fppowtf32.vhdl:3905:33  */
  assign n689 = ~n688;
  /* fppowtf32.vhdl:3905:31  */
  assign n691 = {1'b1, n689};
  /* fppowtf32.vhdl:3906:4  */
  intadder_24_freq500_uid22 additer2_1 (
    .clk(clk),
    .x(eiypb1),
    .y(pp1),
    .cin(n692),
    .r(additer2_1_n693));
  /* fppowtf32.vhdl:3913:26  */
  assign n696 = zfinal_d2[23:9]; // extract
  /* fppowtf32.vhdl:3913:54  */
  assign n697 = dorr_d2 ? n696 : n699;
  /* fppowtf32.vhdl:3914:48  */
  assign n699 = {small_absz0_normd_d1, 4'b0000};
  /* fppowtf32.vhdl:3915:26  */
  assign n700 = {15'b0, squarerin};  //  uext
  /* fppowtf32.vhdl:3915:26  */
  assign n701 = {15'b0, squarerin};  //  uext
  /* fppowtf32.vhdl:3915:26  */
  assign n702 = n700 * n701; // umul
  /* fppowtf32.vhdl:3917:35  */
  assign n703 = z2o2_full_dummy[29:18]; // extract
  /* fppowtf32.vhdl:3918:50  */
  assign n704 = ~z2o2_normal;
  /* fppowtf32.vhdl:3918:48  */
  assign n706 = {12'b111111111111, n704};
  /* fppowtf32.vhdl:3919:4  */
  intadder_24_freq500_uid25 addfinallog1p_normaladder (
    .clk(clk),
    .x(zfinal),
    .y(addfinallog1py),
    .cin(n707),
    .r(addfinallog1p_normaladder_n708));
  /* fppowtf32.vhdl:3927:4  */
  logtable0_freq500_uid27 logtable0 (
    .x(a0),
    .y(logtable0_n711));
  /* fppowtf32.vhdl:3932:4  */
  logtable1_freq500_uid30 logtable1 (
    .x(a1),
    .y(logtable1_n714));
  /* fppowtf32.vhdl:3936:36  */
  assign n718 = {6'b000000, l1};
  /* fppowtf32.vhdl:3937:4  */
  intadder_35_freq500_uid34 adders1 (
    .clk(clk),
    .x(s1),
    .y(sopx1),
    .cin(n719),
    .r(adders1_n720));
  /* fppowtf32.vhdl:3944:62  */
  assign n724 = {11'b00000000000, log1p_normal};
  /* fppowtf32.vhdl:3945:4  */
  intadder_35_freq500_uid37 adderlogf_normal (
    .clk(clk),
    .x(almostlog),
    .y(adderlogf_normaly),
    .cin(n725),
    .r(adderlogf_normal_n726));
  /* fppowtf32.vhdl:3951:4  */
  fixrealkcm_freq500_uid39 mullog2 (
    .clk(clk),
    .x(abse),
    .r(mullog2_n729));
  /* fppowtf32.vhdl:3955:31  */
  assign n733 = {abselog2, 11'b00000000000};
  /* fppowtf32.vhdl:3956:53  */
  assign n734 = logf_normal[34]; // extract
  /* fppowtf32.vhdl:3956:53  */
  assign n735 = logf_normal[34]; // extract
  /* fppowtf32.vhdl:3956:53  */
  assign n736 = logf_normal[34]; // extract
  /* fppowtf32.vhdl:3956:53  */
  assign n737 = logf_normal[34]; // extract
  /* fppowtf32.vhdl:3956:53  */
  assign n738 = logf_normal[34]; // extract
  /* fppowtf32.vhdl:3956:53  */
  assign n739 = logf_normal[34]; // extract
  /* fppowtf32.vhdl:3956:53  */
  assign n740 = logf_normal[34]; // extract
  /* fppowtf32.vhdl:3956:53  */
  assign n741 = logf_normal[34]; // extract
  assign n742 = {n741, n740, n739, n738};
  assign n743 = {n737, n736, n735, n734};
  assign n744 = {n742, n743};
  /* fppowtf32.vhdl:3956:70  */
  assign n745 = {n744, logf_normal};
  /* fppowtf32.vhdl:3958:40  */
  assign n746 = ~sr_d6;
  /* fppowtf32.vhdl:3958:30  */
  assign n747 = n746 ? logf_normal_pad : n748;
  /* fppowtf32.vhdl:3958:50  */
  assign n748 = ~logf_normal_pad;
  /* fppowtf32.vhdl:3959:4  */
  intadder_43_freq500_uid51 lnadder (
    .clk(clk),
    .x(lnaddx),
    .y(lnaddy),
    .cin(sr),
    .r(lnadder_n749));
  /* fppowtf32.vhdl:3965:4  */
  normalizer_z_43_35_18_freq500_uid53 final_norm (
    .clk(clk),
    .x(log_normal),
    .count(final_norm_n752),
    .r(final_norm_n753));
  /* fppowtf32.vhdl:3970:36  */
  assign n758 = z2o2_full_dummy[29:15]; // extract
  /* fppowtf32.vhdl:3971:4  */
  rightshifter15_by_max_14_freq500_uid55 ao_rshift (
    .clk(clk),
    .x(z2o2_small_bs),
    .s(shiftvalinr),
    .r(ao_rshift_n759));
  /* fppowtf32.vhdl:3977:61  */
  assign n762 = z2o2_small_s[28:14]; // extract
  /* fppowtf32.vhdl:3977:47  */
  assign n764 = {11'b00000000000, n762};
  /* fppowtf32.vhdl:3979:33  */
  assign n766 = {small_absz0_normd, 15'b000000000000000};
  /* fppowtf32.vhdl:3980:29  */
  assign n767 = sr_d6 ? z2o2_small : n768;
  /* fppowtf32.vhdl:3980:49  */
  assign n768 = ~z2o2_small;
  /* fppowtf32.vhdl:3981:14  */
  assign n769 = ~sr;
  /* fppowtf32.vhdl:3982:4  */
  intadder_26_freq500_uid57 log_small_adder (
    .clk(clk),
    .x(z_small),
    .y(log_smally),
    .cin(nsrcin),
    .r(log_small_adder_n770));
  /* fppowtf32.vhdl:3989:35  */
  assign n774 = log_small[25]; // extract
  /* fppowtf32.vhdl:3989:21  */
  assign n775 = n774 ? 2'b11 : n780;
  /* fppowtf32.vhdl:3990:35  */
  assign n777 = log_small[25:24]; // extract
  /* fppowtf32.vhdl:3990:56  */
  assign n779 = n777 == 2'b01;
  /* fppowtf32.vhdl:3990:11  */
  assign n780 = n779 ? 2'b10 : 2'b01;
  /* fppowtf32.vhdl:3996:46  */
  assign n784 = {6'b011111, e0_sub};
  /* fppowtf32.vhdl:3996:84  */
  assign n786 = {3'b000, lzo_d3};
  /* fppowtf32.vhdl:3996:57  */
  assign n787 = n784 - n786;
  /* fppowtf32.vhdl:3997:32  */
  assign n788 = log_small[25:2]; // extract
  /* fppowtf32.vhdl:3997:64  */
  assign n789 = log_small[25]; // extract
  /* fppowtf32.vhdl:3997:50  */
  assign n790 = n789 ? n788 : n793;
  /* fppowtf32.vhdl:3998:26  */
  assign n791 = log_small[24:1]; // extract
  /* fppowtf32.vhdl:3998:57  */
  assign n792 = log_small[24]; // extract
  /* fppowtf32.vhdl:3998:12  */
  assign n793 = n792 ? n791 : n794;
  /* fppowtf32.vhdl:3999:26  */
  assign n794 = log_small[23:0]; // extract
  /* fppowtf32.vhdl:4001:33  */
  assign n796 = small_d6 ? e_small_d4 : n799;
  /* fppowtf32.vhdl:4002:48  */
  assign n798 = {3'b000, e_normal};
  /* fppowtf32.vhdl:4002:25  */
  assign n799 = e0offset_d10 - n798;
  /* fppowtf32.vhdl:4003:32  */
  assign n800 = log_small_normd_d5[22:0]; // extract
  /* fppowtf32.vhdl:4003:50  */
  assign n802 = {n800, 1'b0};
  /* fppowtf32.vhdl:4003:56  */
  assign n803 = small_d7 ? n802 : n804;
  /* fppowtf32.vhdl:4004:28  */
  assign n804 = log_normal_normd[33:10]; // extract
  /* fppowtf32.vhdl:4005:18  */
  assign n805 = log_g[3]; // extract
  /* fppowtf32.vhdl:4007:26  */
  assign n806 = log_g[23:4]; // extract
  /* fppowtf32.vhdl:4007:19  */
  assign n807 = {er_d1, n806};
  /* fppowtf32.vhdl:4008:39  */
  assign n809 = {27'b000000000000000000000000000, round};
  /* fppowtf32.vhdl:4009:4  */
  intadder_28_freq500_uid60 finalroundadder (
    .clk(clk),
    .x(frax),
    .y(fray),
    .cin(n810),
    .r(finalroundadder_n811));
  /* fppowtf32.vhdl:4015:36  */
  assign n815 = xexnsgn_d11[2]; // extract
  /* fppowtf32.vhdl:4015:56  */
  assign n816 = xexnsgn_d11[1]; // extract
  /* fppowtf32.vhdl:4015:74  */
  assign n817 = xexnsgn_d11[0]; // extract
  /* fppowtf32.vhdl:4015:60  */
  assign n818 = n816 | n817;
  /* fppowtf32.vhdl:4015:40  */
  assign n819 = n815 & n818;
  /* fppowtf32.vhdl:4015:95  */
  assign n820 = xexnsgn_d11[1]; // extract
  /* fppowtf32.vhdl:4015:114  */
  assign n821 = xexnsgn_d11[0]; // extract
  /* fppowtf32.vhdl:4015:99  */
  assign n822 = n820 & n821;
  /* fppowtf32.vhdl:4015:80  */
  assign n823 = n819 | n822;
  /* fppowtf32.vhdl:4015:18  */
  assign n824 = n823 ? 3'b110 : n829;
  /* fppowtf32.vhdl:4016:53  */
  assign n826 = xexnsgn_d11[2:1]; // extract
  /* fppowtf32.vhdl:4016:66  */
  assign n828 = n826 == 2'b00;
  /* fppowtf32.vhdl:4015:126  */
  assign n829 = n828 ? 3'b101 : n834;
  /* fppowtf32.vhdl:4017:53  */
  assign n831 = xexnsgn_d11[2:1]; // extract
  /* fppowtf32.vhdl:4017:66  */
  assign n833 = n831 == 2'b10;
  /* fppowtf32.vhdl:4016:74  */
  assign n834 = n833 ? 3'b100 : n847;
  /* fppowtf32.vhdl:4018:36  */
  assign n836 = {2'b00, sr_d11};
  /* fppowtf32.vhdl:4018:69  */
  assign n837 = log_normal_normd[34]; // extract
  /* fppowtf32.vhdl:4018:83  */
  assign n838 = ~n837;
  /* fppowtf32.vhdl:4018:102  */
  assign n839 = ~small_d7;
  /* fppowtf32.vhdl:4018:89  */
  assign n840 = n839 & n838;
  /* fppowtf32.vhdl:4018:134  */
  assign n841 = log_small_normd_d5[23]; // extract
  /* fppowtf32.vhdl:4018:142  */
  assign n842 = ~n841;
  /* fppowtf32.vhdl:4018:148  */
  assign n843 = small_d7 & n842;
  /* fppowtf32.vhdl:4018:109  */
  assign n844 = n840 | n843;
  /* fppowtf32.vhdl:4018:187  */
  assign n845 = small_d7 & ufl_d11;
  /* fppowtf32.vhdl:4018:169  */
  assign n846 = n844 | n845;
  /* fppowtf32.vhdl:4017:74  */
  assign n847 = n846 ? n836 : n849;
  /* fppowtf32.vhdl:4019:37  */
  assign n849 = {2'b01, sr_d11};
  /* fppowtf32.vhdl:4020:14  */
  assign n850 = {rexn, efr};
  /* fppowtf32.vhdl:3768:10  */
  always @(posedge clk)
    n851 <= xexnsgn;
  /* fppowtf32.vhdl:3768:10  */
  always @(posedge clk)
    n852 <= xexnsgn_d1;
  /* fppowtf32.vhdl:3768:10  */
  always @(posedge clk)
    n853 <= xexnsgn_d2;
  /* fppowtf32.vhdl:3768:10  */
  always @(posedge clk)
    n854 <= xexnsgn_d3;
  /* fppowtf32.vhdl:3768:10  */
  always @(posedge clk)
    n855 <= xexnsgn_d4;
  /* fppowtf32.vhdl:3768:10  */
  always @(posedge clk)
    n856 <= xexnsgn_d5;
  /* fppowtf32.vhdl:3768:10  */
  always @(posedge clk)
    n857 <= xexnsgn_d6;
  /* fppowtf32.vhdl:3768:10  */
  always @(posedge clk)
    n858 <= xexnsgn_d7;
  /* fppowtf32.vhdl:3768:10  */
  always @(posedge clk)
    n859 <= xexnsgn_d8;
  /* fppowtf32.vhdl:3768:10  */
  always @(posedge clk)
    n860 <= xexnsgn_d9;
  /* fppowtf32.vhdl:3768:10  */
  always @(posedge clk)
    n861 <= xexnsgn_d10;
  /* fppowtf32.vhdl:3768:10  */
  always @(posedge clk)
    n862 <= y0;
  /* fppowtf32.vhdl:3768:10  */
  always @(posedge clk)
    n863 <= sr;
  /* fppowtf32.vhdl:3768:10  */
  always @(posedge clk)
    n864 <= sr_d1;
  /* fppowtf32.vhdl:3768:10  */
  always @(posedge clk)
    n865 <= sr_d2;
  /* fppowtf32.vhdl:3768:10  */
  always @(posedge clk)
    n866 <= sr_d3;
  /* fppowtf32.vhdl:3768:10  */
  always @(posedge clk)
    n867 <= sr_d4;
  /* fppowtf32.vhdl:3768:10  */
  always @(posedge clk)
    n868 <= sr_d5;
  /* fppowtf32.vhdl:3768:10  */
  always @(posedge clk)
    n869 <= sr_d6;
  /* fppowtf32.vhdl:3768:10  */
  always @(posedge clk)
    n870 <= sr_d7;
  /* fppowtf32.vhdl:3768:10  */
  always @(posedge clk)
    n871 <= sr_d8;
  /* fppowtf32.vhdl:3768:10  */
  always @(posedge clk)
    n872 <= sr_d9;
  /* fppowtf32.vhdl:3768:10  */
  always @(posedge clk)
    n873 <= sr_d10;
  /* fppowtf32.vhdl:3768:10  */
  always @(posedge clk)
    n874 <= eeqzero;
  /* fppowtf32.vhdl:3768:10  */
  always @(posedge clk)
    n875 <= eeqzero_d1;
  /* fppowtf32.vhdl:3768:10  */
  always @(posedge clk)
    n876 <= eeqzero_d2;
  /* fppowtf32.vhdl:3768:10  */
  always @(posedge clk)
    n877 <= eeqzero_d3;
  /* fppowtf32.vhdl:3768:10  */
  always @(posedge clk)
    n878 <= lzo;
  /* fppowtf32.vhdl:3768:10  */
  always @(posedge clk)
    n879 <= lzo_d1;
  /* fppowtf32.vhdl:3768:10  */
  always @(posedge clk)
    n880 <= lzo_d2;
  /* fppowtf32.vhdl:3768:10  */
  always @(posedge clk)
    n881 <= pfinal_s;
  /* fppowtf32.vhdl:3768:10  */
  always @(posedge clk)
    n882 <= pfinal_s_d1;
  /* fppowtf32.vhdl:3768:10  */
  always @(posedge clk)
    n883 <= pfinal_s_d2;
  /* fppowtf32.vhdl:3768:10  */
  always @(posedge clk)
    n884 <= dorr;
  /* fppowtf32.vhdl:3768:10  */
  always @(posedge clk)
    n885 <= dorr_d1;
  /* fppowtf32.vhdl:3768:10  */
  always @(posedge clk)
    n886 <= \small ;
  /* fppowtf32.vhdl:3768:10  */
  always @(posedge clk)
    n887 <= small_d1;
  /* fppowtf32.vhdl:3768:10  */
  always @(posedge clk)
    n888 <= small_d2;
  /* fppowtf32.vhdl:3768:10  */
  always @(posedge clk)
    n889 <= small_d3;
  /* fppowtf32.vhdl:3768:10  */
  always @(posedge clk)
    n890 <= small_d4;
  /* fppowtf32.vhdl:3768:10  */
  always @(posedge clk)
    n891 <= small_d5;
  /* fppowtf32.vhdl:3768:10  */
  always @(posedge clk)
    n892 <= small_d6;
  /* fppowtf32.vhdl:3768:10  */
  always @(posedge clk)
    n893 <= small_absz0_normd;
  /* fppowtf32.vhdl:3768:10  */
  always @(posedge clk)
    n894 <= inva0;
  /* fppowtf32.vhdl:3768:10  */
  always @(posedge clk)
    n895 <= a1;
  /* fppowtf32.vhdl:3768:10  */
  always @(posedge clk)
    n896 <= zm1;
  /* fppowtf32.vhdl:3768:10  */
  always @(posedge clk)
    n897 <= zfinal;
  /* fppowtf32.vhdl:3768:10  */
  always @(posedge clk)
    n898 <= zfinal_d1;
  /* fppowtf32.vhdl:3768:10  */
  always @(posedge clk)
    n899 <= ufl;
  /* fppowtf32.vhdl:3768:10  */
  always @(posedge clk)
    n900 <= ufl_d1;
  /* fppowtf32.vhdl:3768:10  */
  always @(posedge clk)
    n901 <= ufl_d2;
  /* fppowtf32.vhdl:3768:10  */
  always @(posedge clk)
    n902 <= ufl_d3;
  /* fppowtf32.vhdl:3768:10  */
  always @(posedge clk)
    n903 <= ufl_d4;
  /* fppowtf32.vhdl:3768:10  */
  always @(posedge clk)
    n904 <= ufl_d5;
  /* fppowtf32.vhdl:3768:10  */
  always @(posedge clk)
    n905 <= ufl_d6;
  /* fppowtf32.vhdl:3768:10  */
  always @(posedge clk)
    n906 <= ufl_d7;
  /* fppowtf32.vhdl:3768:10  */
  always @(posedge clk)
    n907 <= ufl_d8;
  /* fppowtf32.vhdl:3768:10  */
  always @(posedge clk)
    n908 <= ufl_d9;
  /* fppowtf32.vhdl:3768:10  */
  always @(posedge clk)
    n909 <= ufl_d10;
  /* fppowtf32.vhdl:3768:10  */
  always @(posedge clk)
    n910 <= e_small;
  /* fppowtf32.vhdl:3768:10  */
  always @(posedge clk)
    n911 <= e_small_d1;
  /* fppowtf32.vhdl:3768:10  */
  always @(posedge clk)
    n912 <= e_small_d2;
  /* fppowtf32.vhdl:3768:10  */
  always @(posedge clk)
    n913 <= e_small_d3;
  /* fppowtf32.vhdl:3768:10  */
  always @(posedge clk)
    n914 <= log_small_normd;
  /* fppowtf32.vhdl:3768:10  */
  always @(posedge clk)
    n915 <= log_small_normd_d1;
  /* fppowtf32.vhdl:3768:10  */
  always @(posedge clk)
    n916 <= log_small_normd_d2;
  /* fppowtf32.vhdl:3768:10  */
  always @(posedge clk)
    n917 <= log_small_normd_d3;
  /* fppowtf32.vhdl:3768:10  */
  always @(posedge clk)
    n918 <= log_small_normd_d4;
  /* fppowtf32.vhdl:3768:10  */
  always @(posedge clk)
    n919 <= e0offset;
  /* fppowtf32.vhdl:3768:10  */
  always @(posedge clk)
    n920 <= e0offset_d1;
  /* fppowtf32.vhdl:3768:10  */
  always @(posedge clk)
    n921 <= e0offset_d2;
  /* fppowtf32.vhdl:3768:10  */
  always @(posedge clk)
    n922 <= e0offset_d3;
  /* fppowtf32.vhdl:3768:10  */
  always @(posedge clk)
    n923 <= e0offset_d4;
  /* fppowtf32.vhdl:3768:10  */
  always @(posedge clk)
    n924 <= e0offset_d5;
  /* fppowtf32.vhdl:3768:10  */
  always @(posedge clk)
    n925 <= e0offset_d6;
  /* fppowtf32.vhdl:3768:10  */
  always @(posedge clk)
    n926 <= e0offset_d7;
  /* fppowtf32.vhdl:3768:10  */
  always @(posedge clk)
    n927 <= e0offset_d8;
  /* fppowtf32.vhdl:3768:10  */
  always @(posedge clk)
    n928 <= e0offset_d9;
  /* fppowtf32.vhdl:3768:10  */
  always @(posedge clk)
    n929 <= er;
endmodule

module lzc_10_freq500_uid7
  (input  clk,
   input  [9:0] i,
   output [3:0] o);
  wire [14:0] level4;
  wire digit3;
  wire [6:0] level3;
  wire [6:0] level3_d1;
  wire digit2;
  wire digit2_d1;
  wire [2:0] level2;
  wire [1:0] lowbits;
  wire [1:0] outhighbits;
  wire [1:0] outhighbits_d1;
  wire [14:0] n478;
  wire [7:0] n480;
  wire n482;
  wire n483;
  wire [6:0] n485;
  wire [6:0] n486;
  wire [6:0] n487;
  wire [3:0] n489;
  wire n491;
  wire n492;
  wire [2:0] n494;
  wire [2:0] n495;
  wire [2:0] n496;
  wire n499;
  wire n502;
  wire n505;
  wire n508;
  wire [3:0] n510;
  reg [1:0] n511;
  wire [1:0] n512;
  wire [3:0] n514;
  reg [6:0] n515;
  reg n516;
  reg [1:0] n517;
  assign o = n514; //(module output)
  /* fppowtf32.vhdl:2266:8  */
  assign level4 = n478; // (signal)
  /* fppowtf32.vhdl:2268:8  */
  assign digit3 = n483; // (signal)
  /* fppowtf32.vhdl:2270:8  */
  assign level3 = n486; // (signal)
  /* fppowtf32.vhdl:2270:16  */
  assign level3_d1 = n515; // (signal)
  /* fppowtf32.vhdl:2272:8  */
  assign digit2 = n492; // (signal)
  /* fppowtf32.vhdl:2272:16  */
  assign digit2_d1 = n516; // (signal)
  /* fppowtf32.vhdl:2274:8  */
  assign level2 = n495; // (signal)
  /* fppowtf32.vhdl:2276:8  */
  assign lowbits = n511; // (signal)
  /* fppowtf32.vhdl:2278:8  */
  assign outhighbits = n512; // (signal)
  /* fppowtf32.vhdl:2278:21  */
  assign outhighbits_d1 = n517; // (signal)
  /* fppowtf32.vhdl:2290:16  */
  assign n478 = {i, 5'b11111};
  /* fppowtf32.vhdl:2292:28  */
  assign n480 = level4[14:7]; // extract
  /* fppowtf32.vhdl:2292:42  */
  assign n482 = n480 == 8'b00000000;
  /* fppowtf32.vhdl:2292:17  */
  assign n483 = n482 ? 1'b1 : 1'b0;
  /* fppowtf32.vhdl:2293:19  */
  assign n485 = level4[6:0]; // extract
  /* fppowtf32.vhdl:2293:32  */
  assign n486 = digit3 ? n485 : n487;
  /* fppowtf32.vhdl:2293:59  */
  assign n487 = level4[14:8]; // extract
  /* fppowtf32.vhdl:2294:28  */
  assign n489 = level3[6:3]; // extract
  /* fppowtf32.vhdl:2294:41  */
  assign n491 = n489 == 4'b0000;
  /* fppowtf32.vhdl:2294:17  */
  assign n492 = n491 ? 1'b1 : 1'b0;
  /* fppowtf32.vhdl:2295:22  */
  assign n494 = level3_d1[2:0]; // extract
  /* fppowtf32.vhdl:2295:35  */
  assign n495 = digit2_d1 ? n494 : n496;
  /* fppowtf32.vhdl:2295:68  */
  assign n496 = level3_d1[6:4]; // extract
  /* fppowtf32.vhdl:2298:12  */
  assign n499 = level2 == 3'b000;
  /* fppowtf32.vhdl:2299:12  */
  assign n502 = level2 == 3'b001;
  /* fppowtf32.vhdl:2300:12  */
  assign n505 = level2 == 3'b010;
  /* fppowtf32.vhdl:2301:12  */
  assign n508 = level2 == 3'b011;
  assign n510 = {n508, n505, n502, n499};
  /* fppowtf32.vhdl:2297:4  */
  always @*
    case (n510)
      4'b1000: n511 = 2'b01;
      4'b0100: n511 = 2'b01;
      4'b0010: n511 = 2'b10;
      4'b0001: n511 = 2'b11;
      default: n511 = 2'b00;
    endcase
  /* fppowtf32.vhdl:2303:35  */
  assign n512 = {digit3, digit2};
  /* fppowtf32.vhdl:2304:24  */
  assign n514 = {outhighbits_d1, lowbits};
  /* fppowtf32.vhdl:2283:10  */
  always @(posedge clk)
    n515 <= level3;
  /* fppowtf32.vhdl:2283:10  */
  always @(posedge clk)
    n516 <= digit2;
  /* fppowtf32.vhdl:2283:10  */
  always @(posedge clk)
    n517 <= outhighbits;
endmodule

module intadder_19_freq500_uid5
  (input  clk,
   input  [18:0] x,
   input  [18:0] y,
   input  cin,
   output [18:0] r);
  wire [18:0] rtmp;
  wire [18:0] n466;
  wire [18:0] n467;
  wire [18:0] n468;
  assign r = rtmp; //(module output)
  /* fppowtf32.vhdl:2229:8  */
  assign rtmp = n468; // (signal)
  /* fppowtf32.vhdl:2232:14  */
  assign n466 = x + y;
  /* fppowtf32.vhdl:2232:18  */
  assign n467 = {18'b0, cin};  //  uext
  /* fppowtf32.vhdl:2232:18  */
  assign n468 = n466 + n467;
endmodule

module top_module
  (input  clk,
   input  [20:0] X,
   input  [20:0] Y,
   output [20:0] R);
  wire [1:0] flagsx;
  wire signx;
  wire signx_d1;
  wire signx_d2;
  wire [7:0] expfieldx;
  wire [9:0] fracx;
  wire [1:0] flagsy;
  wire signy;
  wire signy_d1;
  wire signy_d2;
  wire signy_d3;
  wire [7:0] expfieldy;
  wire [9:0] fracy;
  wire zerox;
  wire zerox_d1;
  wire zerox_d2;
  wire zerox_d3;
  wire zeroy;
  wire zeroy_d1;
  wire zeroy_d2;
  wire normalx;
  wire normalx_d1;
  wire normalx_d2;
  wire normaly;
  wire normaly_d1;
  wire normaly_d2;
  wire normaly_d3;
  wire infx;
  wire infx_d1;
  wire infx_d2;
  wire infx_d3;
  wire infy;
  wire infy_d1;
  wire infy_d2;
  wire infy_d3;
  wire s_nan_in;
  wire s_nan_in_d1;
  wire s_nan_in_d2;
  wire [17:0] oneexpfrac;
  wire [18:0] expfracx;
  wire [18:0] oneexpfraccompl;
  wire [18:0] cmpxoneres;
  wire xisoneandnormal;
  wire absxgtoneandnormal;
  wire absxgtoneandnormal_d1;
  wire absxgtoneandnormal_d2;
  wire absxgtoneandnormal_d3;
  wire absxltoneandnormal;
  wire absxltoneandnormal_d1;
  wire absxltoneandnormal_d2;
  wire absxltoneandnormal_d3;
  wire [9:0] fracyreverted;
  wire [3:0] z_righty;
  wire [3:0] z_righty_d1;
  wire [8:0] weightlsbypre;
  wire [8:0] weightlsbypre_d1;
  wire [8:0] weightlsbypre_d2;
  wire [8:0] weightlsby;
  wire oddinty;
  wire oddinty_d1;
  wire eveninty;
  wire eveninty_d1;
  wire notintnormaly;
  wire risinfspecialcase;
  wire risinfspecialcase_d1;
  wire risinfspecialcase_d2;
  wire risinfspecialcase_d3;
  wire risinfspecialcase_d4;
  wire risinfspecialcase_d5;
  wire risinfspecialcase_d6;
  wire risinfspecialcase_d7;
  wire risinfspecialcase_d8;
  wire risinfspecialcase_d9;
  wire risinfspecialcase_d10;
  wire risinfspecialcase_d11;
  wire risinfspecialcase_d12;
  wire risinfspecialcase_d13;
  wire risinfspecialcase_d14;
  wire risinfspecialcase_d15;
  wire risinfspecialcase_d16;
  wire risinfspecialcase_d17;
  wire risinfspecialcase_d18;
  wire riszerospecialcase;
  wire riszerospecialcase_d1;
  wire riszerospecialcase_d2;
  wire riszerospecialcase_d3;
  wire riszerospecialcase_d4;
  wire riszerospecialcase_d5;
  wire riszerospecialcase_d6;
  wire riszerospecialcase_d7;
  wire riszerospecialcase_d8;
  wire riszerospecialcase_d9;
  wire riszerospecialcase_d10;
  wire riszerospecialcase_d11;
  wire riszerospecialcase_d12;
  wire riszerospecialcase_d13;
  wire riszerospecialcase_d14;
  wire riszerospecialcase_d15;
  wire riszerospecialcase_d16;
  wire riszerospecialcase_d17;
  wire riszerospecialcase_d18;
  wire risone;
  wire risone_d1;
  wire risone_d2;
  wire risone_d3;
  wire risone_d4;
  wire risone_d5;
  wire risone_d6;
  wire risone_d7;
  wire risone_d8;
  wire risone_d9;
  wire risone_d10;
  wire risone_d11;
  wire risone_d12;
  wire risone_d13;
  wire risone_d14;
  wire risone_d15;
  wire risone_d16;
  wire risone_d17;
  wire risone_d18;
  wire risone_d19;
  wire risone_d20;
  wire risone_d21;
  wire risnan;
  wire risnan_d1;
  wire risnan_d2;
  wire risnan_d3;
  wire risnan_d4;
  wire risnan_d5;
  wire risnan_d6;
  wire risnan_d7;
  wire risnan_d8;
  wire risnan_d9;
  wire risnan_d10;
  wire risnan_d11;
  wire risnan_d12;
  wire risnan_d13;
  wire risnan_d14;
  wire risnan_d15;
  wire risnan_d16;
  wire risnan_d17;
  wire risnan_d18;
  wire risnan_d19;
  wire signr;
  wire signr_d1;
  wire signr_d2;
  wire signr_d3;
  wire signr_d4;
  wire signr_d5;
  wire signr_d6;
  wire signr_d7;
  wire signr_d8;
  wire signr_d9;
  wire signr_d10;
  wire signr_d11;
  wire signr_d12;
  wire signr_d13;
  wire signr_d14;
  wire signr_d15;
  wire signr_d16;
  wire signr_d17;
  wire signr_d18;
  wire signr_d19;
  wire [30:0] login;
  wire [30:0] lnx;
  wire [31:0] p;
  wire [20:0] e;
  wire [20:0] e_d1;
  wire [1:0] flagse;
  wire [1:0] flagse_d1;
  wire riszerofromexp;
  wire riszero;
  wire risinffromexp;
  wire risinf;
  wire [1:0] flagr;
  wire [17:0] r_expfrac;
  wire [1:0] n136;
  wire n137;
  wire [7:0] n138;
  wire [9:0] n139;
  wire [1:0] n140;
  wire n141;
  wire [7:0] n142;
  wire [9:0] n143;
  wire n146;
  wire n147;
  wire n151;
  wire n152;
  wire n156;
  wire n157;
  wire n161;
  wire n162;
  wire n166;
  wire n167;
  wire n171;
  wire n172;
  wire n176;
  wire n178;
  wire n179;
  wire n180;
  wire [8:0] n184;
  wire [18:0] n185;
  wire [17:0] n186;
  wire [18:0] n188;
  localparam n189 = 1'b1;
  wire [18:0] cmpxone_n190;
  wire [20:0] n195;
  wire n196;
  wire n197;
  wire n199;
  wire n200;
  wire n201;
  wire n202;
  wire n203;
  wire n204;
  wire n205;
  wire n206;
  wire n207;
  wire [1:0] n208;
  wire n209;
  wire [2:0] n210;
  wire n211;
  wire [3:0] n212;
  wire n213;
  wire [4:0] n214;
  wire n215;
  wire [5:0] n216;
  wire n217;
  wire [6:0] n218;
  wire n219;
  wire [7:0] n220;
  wire n221;
  wire [8:0] n222;
  wire n223;
  wire [9:0] n224;
  wire [3:0] fppow_8_10_freq500_uid2right1counter_n225;
  wire [8:0] n229;
  wire [8:0] n231;
  wire [8:0] n232;
  wire [8:0] n233;
  wire n235;
  wire n236;
  wire n238;
  wire n239;
  wire n240;
  wire n241;
  wire n242;
  wire n244;
  wire n245;
  wire n247;
  wire n248;
  wire n249;
  wire n250;
  wire n251;
  wire n252;
  wire n253;
  wire n254;
  wire n255;
  wire n256;
  wire n257;
  wire n258;
  wire n259;
  wire n260;
  wire n261;
  wire n262;
  wire n263;
  wire n264;
  wire n265;
  wire n266;
  wire n267;
  wire n268;
  wire n269;
  wire n270;
  wire n271;
  wire n272;
  wire n273;
  wire n274;
  wire n275;
  wire n276;
  wire n277;
  wire n278;
  wire n279;
  wire n280;
  wire n281;
  wire n282;
  wire n283;
  wire n284;
  wire n285;
  wire n286;
  wire n287;
  wire n288;
  wire n289;
  wire n290;
  wire n291;
  wire n292;
  wire n293;
  wire [2:0] n295;
  wire [10:0] n296;
  wire [20:0] n297;
  wire [30:0] n299;
  wire [30:0] fppow_8_10_freq500_uid2log_n300;
  wire [31:0] fppow_8_10_freq500_uid2mult_n303;
  wire [20:0] fppow_8_10_freq500_uid2exp_n306;
  wire [1:0] n309;
  wire n312;
  wire n313;
  wire n315;
  wire n318;
  wire n319;
  wire n321;
  wire [1:0] n323;
  wire [1:0] n325;
  wire [1:0] n327;
  wire [17:0] n330;
  wire [17:0] n331;
  wire [2:0] n332;
  wire [20:0] n333;
  reg n334;
  reg n335;
  reg n336;
  reg n337;
  reg n338;
  reg n339;
  reg n340;
  reg n341;
  reg n342;
  reg n343;
  reg n344;
  reg n345;
  reg n346;
  reg n347;
  reg n348;
  reg n349;
  reg n350;
  reg n351;
  reg n352;
  reg n353;
  reg n354;
  reg n355;
  reg n356;
  reg n357;
  reg n358;
  reg n359;
  reg n360;
  reg n361;
  reg n362;
  reg [3:0] n363;
  reg [8:0] n364;
  reg [8:0] n365;
  reg n366;
  reg n367;
  reg n368;
  reg n369;
  reg n370;
  reg n371;
  reg n372;
  reg n373;
  reg n374;
  reg n375;
  reg n376;
  reg n377;
  reg n378;
  reg n379;
  reg n380;
  reg n381;
  reg n382;
  reg n383;
  reg n384;
  reg n385;
  reg n386;
  reg n387;
  reg n388;
  reg n389;
  reg n390;
  reg n391;
  reg n392;
  reg n393;
  reg n394;
  reg n395;
  reg n396;
  reg n397;
  reg n398;
  reg n399;
  reg n400;
  reg n401;
  reg n402;
  reg n403;
  reg n404;
  reg n405;
  reg n406;
  reg n407;
  reg n408;
  reg n409;
  reg n410;
  reg n411;
  reg n412;
  reg n413;
  reg n414;
  reg n415;
  reg n416;
  reg n417;
  reg n418;
  reg n419;
  reg n420;
  reg n421;
  reg n422;
  reg n423;
  reg n424;
  reg n425;
  reg n426;
  reg n427;
  reg n428;
  reg n429;
  reg n430;
  reg n431;
  reg n432;
  reg n433;
  reg n434;
  reg n435;
  reg n436;
  reg n437;
  reg n438;
  reg n439;
  reg n440;
  reg n441;
  reg n442;
  reg n443;
  reg n444;
  reg n445;
  reg n446;
  reg n447;
  reg n448;
  reg n449;
  reg n450;
  reg n451;
  reg n452;
  reg n453;
  reg n454;
  reg n455;
  reg n456;
  reg n457;
  reg n458;
  reg n459;
  reg n460;
  reg n461;
  reg n462;
  reg [20:0] n463;
  reg [1:0] n464;
  assign R = n333; //(module output)
  /* fppowtf32.vhdl:5790:8  */
  assign flagsx = n136; // (signal)
  /* fppowtf32.vhdl:5792:8  */
  assign signx = n137; // (signal)
  /* fppowtf32.vhdl:5792:15  */
  assign signx_d1 = n334; // (signal)
  /* fppowtf32.vhdl:5792:25  */
  assign signx_d2 = n335; // (signal)
  /* fppowtf32.vhdl:5794:8  */
  assign expfieldx = n138; // (signal)
  /* fppowtf32.vhdl:5796:8  */
  assign fracx = n139; // (signal)
  /* fppowtf32.vhdl:5798:8  */
  assign flagsy = n140; // (signal)
  /* fppowtf32.vhdl:5800:8  */
  assign signy = n141; // (signal)
  /* fppowtf32.vhdl:5800:15  */
  assign signy_d1 = n336; // (signal)
  /* fppowtf32.vhdl:5800:25  */
  assign signy_d2 = n337; // (signal)
  /* fppowtf32.vhdl:5800:35  */
  assign signy_d3 = n338; // (signal)
  /* fppowtf32.vhdl:5802:8  */
  assign expfieldy = n142; // (signal)
  /* fppowtf32.vhdl:5804:8  */
  assign fracy = n143; // (signal)
  /* fppowtf32.vhdl:5806:8  */
  assign zerox = n147; // (signal)
  /* fppowtf32.vhdl:5806:15  */
  assign zerox_d1 = n339; // (signal)
  /* fppowtf32.vhdl:5806:25  */
  assign zerox_d2 = n340; // (signal)
  /* fppowtf32.vhdl:5806:35  */
  assign zerox_d3 = n341; // (signal)
  /* fppowtf32.vhdl:5808:8  */
  assign zeroy = n152; // (signal)
  /* fppowtf32.vhdl:5808:15  */
  assign zeroy_d1 = n342; // (signal)
  /* fppowtf32.vhdl:5808:25  */
  assign zeroy_d2 = n343; // (signal)
  /* fppowtf32.vhdl:5810:8  */
  assign normalx = n157; // (signal)
  /* fppowtf32.vhdl:5810:17  */
  assign normalx_d1 = n344; // (signal)
  /* fppowtf32.vhdl:5810:29  */
  assign normalx_d2 = n345; // (signal)
  /* fppowtf32.vhdl:5812:8  */
  assign normaly = n162; // (signal)
  /* fppowtf32.vhdl:5812:17  */
  assign normaly_d1 = n346; // (signal)
  /* fppowtf32.vhdl:5812:29  */
  assign normaly_d2 = n347; // (signal)
  /* fppowtf32.vhdl:5812:41  */
  assign normaly_d3 = n348; // (signal)
  /* fppowtf32.vhdl:5814:8  */
  assign infx = n167; // (signal)
  /* fppowtf32.vhdl:5814:14  */
  assign infx_d1 = n349; // (signal)
  /* fppowtf32.vhdl:5814:23  */
  assign infx_d2 = n350; // (signal)
  /* fppowtf32.vhdl:5814:32  */
  assign infx_d3 = n351; // (signal)
  /* fppowtf32.vhdl:5816:8  */
  assign infy = n172; // (signal)
  /* fppowtf32.vhdl:5816:14  */
  assign infy_d1 = n352; // (signal)
  /* fppowtf32.vhdl:5816:23  */
  assign infy_d2 = n353; // (signal)
  /* fppowtf32.vhdl:5816:32  */
  assign infy_d3 = n354; // (signal)
  /* fppowtf32.vhdl:5818:8  */
  assign s_nan_in = n180; // (signal)
  /* fppowtf32.vhdl:5818:18  */
  assign s_nan_in_d1 = n355; // (signal)
  /* fppowtf32.vhdl:5818:31  */
  assign s_nan_in_d2 = n356; // (signal)
  /* fppowtf32.vhdl:5820:8  */
  assign oneexpfrac = 18'b011111110000000000; // (signal)
  /* fppowtf32.vhdl:5822:8  */
  assign expfracx = n185; // (signal)
  /* fppowtf32.vhdl:5824:8  */
  assign oneexpfraccompl = n188; // (signal)
  /* fppowtf32.vhdl:5826:8  */
  assign cmpxoneres = cmpxone_n190; // (signal)
  /* fppowtf32.vhdl:5828:8  */
  assign xisoneandnormal = n197; // (signal)
  /* fppowtf32.vhdl:5830:8  */
  assign absxgtoneandnormal = n203; // (signal)
  /* fppowtf32.vhdl:5830:28  */
  assign absxgtoneandnormal_d1 = n357; // (signal)
  /* fppowtf32.vhdl:5830:51  */
  assign absxgtoneandnormal_d2 = n358; // (signal)
  /* fppowtf32.vhdl:5830:74  */
  assign absxgtoneandnormal_d3 = n359; // (signal)
  /* fppowtf32.vhdl:5832:8  */
  assign absxltoneandnormal = n205; // (signal)
  /* fppowtf32.vhdl:5832:28  */
  assign absxltoneandnormal_d1 = n360; // (signal)
  /* fppowtf32.vhdl:5832:51  */
  assign absxltoneandnormal_d2 = n361; // (signal)
  /* fppowtf32.vhdl:5832:74  */
  assign absxltoneandnormal_d3 = n362; // (signal)
  /* fppowtf32.vhdl:5834:8  */
  assign fracyreverted = n224; // (signal)
  /* fppowtf32.vhdl:5836:8  */
  assign z_righty = fppow_8_10_freq500_uid2right1counter_n225; // (signal)
  /* fppowtf32.vhdl:5836:18  */
  assign z_righty_d1 = n363; // (signal)
  /* fppowtf32.vhdl:5838:8  */
  assign weightlsbypre = n231; // (signal)
  /* fppowtf32.vhdl:5838:23  */
  assign weightlsbypre_d1 = n364; // (signal)
  /* fppowtf32.vhdl:5838:41  */
  assign weightlsbypre_d2 = n365; // (signal)
  /* fppowtf32.vhdl:5840:8  */
  assign weightlsby = n233; // (signal)
  /* fppowtf32.vhdl:5842:8  */
  assign oddinty = n236; // (signal)
  /* fppowtf32.vhdl:5842:17  */
  assign oddinty_d1 = n366; // (signal)
  /* fppowtf32.vhdl:5844:8  */
  assign eveninty = n242; // (signal)
  /* fppowtf32.vhdl:5844:18  */
  assign eveninty_d1 = n367; // (signal)
  /* fppowtf32.vhdl:5846:8  */
  assign notintnormaly = n245; // (signal)
  /* fppowtf32.vhdl:5848:8  */
  assign risinfspecialcase = n263; // (signal)
  /* fppowtf32.vhdl:5848:27  */
  assign risinfspecialcase_d1 = n368; // (signal)
  /* fppowtf32.vhdl:5848:49  */
  assign risinfspecialcase_d2 = n369; // (signal)
  /* fppowtf32.vhdl:5848:71  */
  assign risinfspecialcase_d3 = n370; // (signal)
  /* fppowtf32.vhdl:5848:93  */
  assign risinfspecialcase_d4 = n371; // (signal)
  /* fppowtf32.vhdl:5848:115  */
  assign risinfspecialcase_d5 = n372; // (signal)
  /* fppowtf32.vhdl:5848:137  */
  assign risinfspecialcase_d6 = n373; // (signal)
  /* fppowtf32.vhdl:5848:159  */
  assign risinfspecialcase_d7 = n374; // (signal)
  /* fppowtf32.vhdl:5848:181  */
  assign risinfspecialcase_d8 = n375; // (signal)
  /* fppowtf32.vhdl:5848:203  */
  assign risinfspecialcase_d9 = n376; // (signal)
  /* fppowtf32.vhdl:5848:225  */
  assign risinfspecialcase_d10 = n377; // (signal)
  /* fppowtf32.vhdl:5848:248  */
  assign risinfspecialcase_d11 = n378; // (signal)
  /* fppowtf32.vhdl:5848:271  */
  assign risinfspecialcase_d12 = n379; // (signal)
  /* fppowtf32.vhdl:5848:294  */
  assign risinfspecialcase_d13 = n380; // (signal)
  /* fppowtf32.vhdl:5848:317  */
  assign risinfspecialcase_d14 = n381; // (signal)
  /* fppowtf32.vhdl:5848:340  */
  assign risinfspecialcase_d15 = n382; // (signal)
  /* fppowtf32.vhdl:5848:363  */
  assign risinfspecialcase_d16 = n383; // (signal)
  /* fppowtf32.vhdl:5848:386  */
  assign risinfspecialcase_d17 = n384; // (signal)
  /* fppowtf32.vhdl:5848:409  */
  assign risinfspecialcase_d18 = n385; // (signal)
  /* fppowtf32.vhdl:5850:8  */
  assign riszerospecialcase = n281; // (signal)
  /* fppowtf32.vhdl:5850:28  */
  assign riszerospecialcase_d1 = n386; // (signal)
  /* fppowtf32.vhdl:5850:51  */
  assign riszerospecialcase_d2 = n387; // (signal)
  /* fppowtf32.vhdl:5850:74  */
  assign riszerospecialcase_d3 = n388; // (signal)
  /* fppowtf32.vhdl:5850:97  */
  assign riszerospecialcase_d4 = n389; // (signal)
  /* fppowtf32.vhdl:5850:120  */
  assign riszerospecialcase_d5 = n390; // (signal)
  /* fppowtf32.vhdl:5850:143  */
  assign riszerospecialcase_d6 = n391; // (signal)
  /* fppowtf32.vhdl:5850:166  */
  assign riszerospecialcase_d7 = n392; // (signal)
  /* fppowtf32.vhdl:5850:189  */
  assign riszerospecialcase_d8 = n393; // (signal)
  /* fppowtf32.vhdl:5850:212  */
  assign riszerospecialcase_d9 = n394; // (signal)
  /* fppowtf32.vhdl:5850:235  */
  assign riszerospecialcase_d10 = n395; // (signal)
  /* fppowtf32.vhdl:5850:259  */
  assign riszerospecialcase_d11 = n396; // (signal)
  /* fppowtf32.vhdl:5850:283  */
  assign riszerospecialcase_d12 = n397; // (signal)
  /* fppowtf32.vhdl:5850:307  */
  assign riszerospecialcase_d13 = n398; // (signal)
  /* fppowtf32.vhdl:5850:331  */
  assign riszerospecialcase_d14 = n399; // (signal)
  /* fppowtf32.vhdl:5850:355  */
  assign riszerospecialcase_d15 = n400; // (signal)
  /* fppowtf32.vhdl:5850:379  */
  assign riszerospecialcase_d16 = n401; // (signal)
  /* fppowtf32.vhdl:5850:403  */
  assign riszerospecialcase_d17 = n402; // (signal)
  /* fppowtf32.vhdl:5850:427  */
  assign riszerospecialcase_d18 = n403; // (signal)
  /* fppowtf32.vhdl:5852:8  */
  assign risone = n287; // (signal)
  /* fppowtf32.vhdl:5852:16  */
  assign risone_d1 = n404; // (signal)
  /* fppowtf32.vhdl:5852:27  */
  assign risone_d2 = n405; // (signal)
  /* fppowtf32.vhdl:5852:38  */
  assign risone_d3 = n406; // (signal)
  /* fppowtf32.vhdl:5852:49  */
  assign risone_d4 = n407; // (signal)
  /* fppowtf32.vhdl:5852:60  */
  assign risone_d5 = n408; // (signal)
  /* fppowtf32.vhdl:5852:71  */
  assign risone_d6 = n409; // (signal)
  /* fppowtf32.vhdl:5852:82  */
  assign risone_d7 = n410; // (signal)
  /* fppowtf32.vhdl:5852:93  */
  assign risone_d8 = n411; // (signal)
  /* fppowtf32.vhdl:5852:104  */
  assign risone_d9 = n412; // (signal)
  /* fppowtf32.vhdl:5852:115  */
  assign risone_d10 = n413; // (signal)
  /* fppowtf32.vhdl:5852:127  */
  assign risone_d11 = n414; // (signal)
  /* fppowtf32.vhdl:5852:139  */
  assign risone_d12 = n415; // (signal)
  /* fppowtf32.vhdl:5852:151  */
  assign risone_d13 = n416; // (signal)
  /* fppowtf32.vhdl:5852:163  */
  assign risone_d14 = n417; // (signal)
  /* fppowtf32.vhdl:5852:175  */
  assign risone_d15 = n418; // (signal)
  /* fppowtf32.vhdl:5852:187  */
  assign risone_d16 = n419; // (signal)
  /* fppowtf32.vhdl:5852:199  */
  assign risone_d17 = n420; // (signal)
  /* fppowtf32.vhdl:5852:211  */
  assign risone_d18 = n421; // (signal)
  /* fppowtf32.vhdl:5852:223  */
  assign risone_d19 = n422; // (signal)
  /* fppowtf32.vhdl:5852:235  */
  assign risone_d20 = n423; // (signal)
  /* fppowtf32.vhdl:5852:247  */
  assign risone_d21 = n424; // (signal)
  /* fppowtf32.vhdl:5854:8  */
  assign risnan = n292; // (signal)
  /* fppowtf32.vhdl:5854:16  */
  assign risnan_d1 = n425; // (signal)
  /* fppowtf32.vhdl:5854:27  */
  assign risnan_d2 = n426; // (signal)
  /* fppowtf32.vhdl:5854:38  */
  assign risnan_d3 = n427; // (signal)
  /* fppowtf32.vhdl:5854:49  */
  assign risnan_d4 = n428; // (signal)
  /* fppowtf32.vhdl:5854:60  */
  assign risnan_d5 = n429; // (signal)
  /* fppowtf32.vhdl:5854:71  */
  assign risnan_d6 = n430; // (signal)
  /* fppowtf32.vhdl:5854:82  */
  assign risnan_d7 = n431; // (signal)
  /* fppowtf32.vhdl:5854:93  */
  assign risnan_d8 = n432; // (signal)
  /* fppowtf32.vhdl:5854:104  */
  assign risnan_d9 = n433; // (signal)
  /* fppowtf32.vhdl:5854:115  */
  assign risnan_d10 = n434; // (signal)
  /* fppowtf32.vhdl:5854:127  */
  assign risnan_d11 = n435; // (signal)
  /* fppowtf32.vhdl:5854:139  */
  assign risnan_d12 = n436; // (signal)
  /* fppowtf32.vhdl:5854:151  */
  assign risnan_d13 = n437; // (signal)
  /* fppowtf32.vhdl:5854:163  */
  assign risnan_d14 = n438; // (signal)
  /* fppowtf32.vhdl:5854:175  */
  assign risnan_d15 = n439; // (signal)
  /* fppowtf32.vhdl:5854:187  */
  assign risnan_d16 = n440; // (signal)
  /* fppowtf32.vhdl:5854:199  */
  assign risnan_d17 = n441; // (signal)
  /* fppowtf32.vhdl:5854:211  */
  assign risnan_d18 = n442; // (signal)
  /* fppowtf32.vhdl:5854:223  */
  assign risnan_d19 = n443; // (signal)
  /* fppowtf32.vhdl:5856:8  */
  assign signr = n293; // (signal)
  /* fppowtf32.vhdl:5856:15  */
  assign signr_d1 = n444; // (signal)
  /* fppowtf32.vhdl:5856:25  */
  assign signr_d2 = n445; // (signal)
  /* fppowtf32.vhdl:5856:35  */
  assign signr_d3 = n446; // (signal)
  /* fppowtf32.vhdl:5856:45  */
  assign signr_d4 = n447; // (signal)
  /* fppowtf32.vhdl:5856:55  */
  assign signr_d5 = n448; // (signal)
  /* fppowtf32.vhdl:5856:65  */
  assign signr_d6 = n449; // (signal)
  /* fppowtf32.vhdl:5856:75  */
  assign signr_d7 = n450; // (signal)
  /* fppowtf32.vhdl:5856:85  */
  assign signr_d8 = n451; // (signal)
  /* fppowtf32.vhdl:5856:95  */
  assign signr_d9 = n452; // (signal)
  /* fppowtf32.vhdl:5856:105  */
  assign signr_d10 = n453; // (signal)
  /* fppowtf32.vhdl:5856:116  */
  assign signr_d11 = n454; // (signal)
  /* fppowtf32.vhdl:5856:127  */
  assign signr_d12 = n455; // (signal)
  /* fppowtf32.vhdl:5856:138  */
  assign signr_d13 = n456; // (signal)
  /* fppowtf32.vhdl:5856:149  */
  assign signr_d14 = n457; // (signal)
  /* fppowtf32.vhdl:5856:160  */
  assign signr_d15 = n458; // (signal)
  /* fppowtf32.vhdl:5856:171  */
  assign signr_d16 = n459; // (signal)
  /* fppowtf32.vhdl:5856:182  */
  assign signr_d17 = n460; // (signal)
  /* fppowtf32.vhdl:5856:193  */
  assign signr_d18 = n461; // (signal)
  /* fppowtf32.vhdl:5856:204  */
  assign signr_d19 = n462; // (signal)
  /* fppowtf32.vhdl:5858:8  */
  assign login = n299; // (signal)
  /* fppowtf32.vhdl:5860:8  */
  assign lnx = fppow_8_10_freq500_uid2log_n300; // (signal)
  /* fppowtf32.vhdl:5862:8  */
  assign p = fppow_8_10_freq500_uid2mult_n303; // (signal)
  /* fppowtf32.vhdl:5864:8  */
  assign e = fppow_8_10_freq500_uid2exp_n306; // (signal)
  /* fppowtf32.vhdl:5864:11  */
  assign e_d1 = n463; // (signal)
  /* fppowtf32.vhdl:5866:8  */
  assign flagse = n309; // (signal)
  /* fppowtf32.vhdl:5866:16  */
  assign flagse_d1 = n464; // (signal)
  /* fppowtf32.vhdl:5868:8  */
  assign riszerofromexp = n313; // (signal)
  /* fppowtf32.vhdl:5870:8  */
  assign riszero = n315; // (signal)
  /* fppowtf32.vhdl:5872:8  */
  assign risinffromexp = n319; // (signal)
  /* fppowtf32.vhdl:5874:8  */
  assign risinf = n321; // (signal)
  /* fppowtf32.vhdl:5876:8  */
  assign flagr = n323; // (signal)
  /* fppowtf32.vhdl:5878:8  */
  assign r_expfrac = n330; // (signal)
  /* fppowtf32.vhdl:6019:15  */
  assign n136 = X[20:19]; // extract
  /* fppowtf32.vhdl:6020:14  */
  assign n137 = X[18]; // extract
  /* fppowtf32.vhdl:6021:18  */
  assign n138 = X[17:10]; // extract
  /* fppowtf32.vhdl:6022:14  */
  assign n139 = X[9:0]; // extract
  /* fppowtf32.vhdl:6023:15  */
  assign n140 = Y[20:19]; // extract
  /* fppowtf32.vhdl:6024:14  */
  assign n141 = Y[18]; // extract
  /* fppowtf32.vhdl:6025:18  */
  assign n142 = Y[17:10]; // extract
  /* fppowtf32.vhdl:6026:14  */
  assign n143 = Y[9:0]; // extract
  /* fppowtf32.vhdl:6029:28  */
  assign n146 = flagsx == 2'b00;
  /* fppowtf32.vhdl:6029:17  */
  assign n147 = n146 ? 1'b1 : 1'b0;
  /* fppowtf32.vhdl:6030:28  */
  assign n151 = flagsy == 2'b00;
  /* fppowtf32.vhdl:6030:17  */
  assign n152 = n151 ? 1'b1 : 1'b0;
  /* fppowtf32.vhdl:6032:30  */
  assign n156 = flagsx == 2'b01;
  /* fppowtf32.vhdl:6032:19  */
  assign n157 = n156 ? 1'b1 : 1'b0;
  /* fppowtf32.vhdl:6033:30  */
  assign n161 = flagsy == 2'b01;
  /* fppowtf32.vhdl:6033:19  */
  assign n162 = n161 ? 1'b1 : 1'b0;
  /* fppowtf32.vhdl:6035:27  */
  assign n166 = flagsx == 2'b10;
  /* fppowtf32.vhdl:6035:16  */
  assign n167 = n166 ? 1'b1 : 1'b0;
  /* fppowtf32.vhdl:6036:27  */
  assign n171 = flagsy == 2'b10;
  /* fppowtf32.vhdl:6036:16  */
  assign n172 = n171 ? 1'b1 : 1'b0;
  /* fppowtf32.vhdl:6038:31  */
  assign n176 = flagsx == 2'b11;
  /* fppowtf32.vhdl:6038:46  */
  assign n178 = flagsy == 2'b11;
  /* fppowtf32.vhdl:6038:37  */
  assign n179 = n176 | n178;
  /* fppowtf32.vhdl:6038:20  */
  assign n180 = n179 ? 1'b1 : 1'b0;
  /* fppowtf32.vhdl:6041:19  */
  assign n184 = {1'b0, expfieldx};
  /* fppowtf32.vhdl:6041:31  */
  assign n185 = {n184, fracx};
  /* fppowtf32.vhdl:6042:30  */
  assign n186 = ~oneexpfrac;
  /* fppowtf32.vhdl:6042:27  */
  assign n188 = {1'b1, n186};
  /* fppowtf32.vhdl:6043:4  */
  intadder_19_freq500_uid5 cmpxone (
    .clk(clk),
    .x(expfracx),
    .y(oneexpfraccompl),
    .cin(n189),
    .r(cmpxone_n190));
  /* fppowtf32.vhdl:6049:43  */
  assign n195 = {3'b010, oneexpfrac};
  /* fppowtf32.vhdl:6049:34  */
  assign n196 = X == n195;
  /* fppowtf32.vhdl:6049:27  */
  assign n197 = n196 ? 1'b1 : 1'b0;
  /* fppowtf32.vhdl:6050:39  */
  assign n199 = ~xisoneandnormal;
  /* fppowtf32.vhdl:6050:34  */
  assign n200 = normalx & n199;
  /* fppowtf32.vhdl:6050:79  */
  assign n201 = cmpxoneres[18]; // extract
  /* fppowtf32.vhdl:6050:65  */
  assign n202 = ~n201;
  /* fppowtf32.vhdl:6050:60  */
  assign n203 = n200 & n202;
  /* fppowtf32.vhdl:6051:48  */
  assign n204 = cmpxoneres[18]; // extract
  /* fppowtf32.vhdl:6051:34  */
  assign n205 = normalx & n204;
  /* fppowtf32.vhdl:6052:26  */
  assign n206 = fracy[0]; // extract
  /* fppowtf32.vhdl:6052:35  */
  assign n207 = fracy[1]; // extract
  /* fppowtf32.vhdl:6052:29  */
  assign n208 = {n206, n207};
  /* fppowtf32.vhdl:6052:44  */
  assign n209 = fracy[2]; // extract
  /* fppowtf32.vhdl:6052:38  */
  assign n210 = {n208, n209};
  /* fppowtf32.vhdl:6052:53  */
  assign n211 = fracy[3]; // extract
  /* fppowtf32.vhdl:6052:47  */
  assign n212 = {n210, n211};
  /* fppowtf32.vhdl:6052:62  */
  assign n213 = fracy[4]; // extract
  /* fppowtf32.vhdl:6052:56  */
  assign n214 = {n212, n213};
  /* fppowtf32.vhdl:6052:71  */
  assign n215 = fracy[5]; // extract
  /* fppowtf32.vhdl:6052:65  */
  assign n216 = {n214, n215};
  /* fppowtf32.vhdl:6052:80  */
  assign n217 = fracy[6]; // extract
  /* fppowtf32.vhdl:6052:74  */
  assign n218 = {n216, n217};
  /* fppowtf32.vhdl:6052:89  */
  assign n219 = fracy[7]; // extract
  /* fppowtf32.vhdl:6052:83  */
  assign n220 = {n218, n219};
  /* fppowtf32.vhdl:6052:98  */
  assign n221 = fracy[8]; // extract
  /* fppowtf32.vhdl:6052:92  */
  assign n222 = {n220, n221};
  /* fppowtf32.vhdl:6052:107  */
  assign n223 = fracy[9]; // extract
  /* fppowtf32.vhdl:6052:101  */
  assign n224 = {n222, n223};
  /* fppowtf32.vhdl:6053:4  */
  lzc_10_freq500_uid7 fppow_8_10_freq500_uid2right1counter (
    .clk(clk),
    .i(fracyreverted),
    .o(fppow_8_10_freq500_uid2right1counter_n225));
  /* fppowtf32.vhdl:6058:26  */
  assign n229 = {1'b0, expfieldy};
  /* fppowtf32.vhdl:6058:38  */
  assign n231 = n229 - 9'b010001001;
  /* fppowtf32.vhdl:6059:35  */
  assign n232 = {5'b0, z_righty_d1};  //  uext
  /* fppowtf32.vhdl:6059:35  */
  assign n233 = weightlsbypre_d2 + n232;
  /* fppowtf32.vhdl:6060:42  */
  assign n235 = weightlsby == 9'b000000000;
  /* fppowtf32.vhdl:6060:26  */
  assign n236 = n235 ? normaly_d2 : 1'b0;
  /* fppowtf32.vhdl:6061:42  */
  assign n238 = weightlsby[8]; // extract
  /* fppowtf32.vhdl:6061:46  */
  assign n239 = ~n238;
  /* fppowtf32.vhdl:6061:62  */
  assign n240 = ~oddinty;
  /* fppowtf32.vhdl:6061:51  */
  assign n241 = n240 & n239;
  /* fppowtf32.vhdl:6061:27  */
  assign n242 = n241 ? normaly_d2 : 1'b0;
  /* fppowtf32.vhdl:6062:47  */
  assign n244 = weightlsby[8]; // extract
  /* fppowtf32.vhdl:6062:32  */
  assign n245 = n244 ? normaly_d2 : 1'b0;
  /* fppowtf32.vhdl:6066:38  */
  assign n247 = oddinty_d1 | eveninty_d1;
  /* fppowtf32.vhdl:6066:21  */
  assign n248 = zerox_d3 & n247;
  /* fppowtf32.vhdl:6066:55  */
  assign n249 = n248 & signy_d3;
  /* fppowtf32.vhdl:6067:20  */
  assign n250 = zerox_d3 & infy_d3;
  /* fppowtf32.vhdl:6067:32  */
  assign n251 = n250 & signy_d3;
  /* fppowtf32.vhdl:6067:7  */
  assign n252 = n249 | n251;
  /* fppowtf32.vhdl:6068:35  */
  assign n253 = absxgtoneandnormal_d3 & infy_d3;
  /* fppowtf32.vhdl:6068:53  */
  assign n254 = ~signy_d3;
  /* fppowtf32.vhdl:6068:49  */
  assign n255 = n253 & n254;
  /* fppowtf32.vhdl:6068:7  */
  assign n256 = n252 | n255;
  /* fppowtf32.vhdl:6069:35  */
  assign n257 = absxltoneandnormal_d3 & infy_d3;
  /* fppowtf32.vhdl:6069:49  */
  assign n258 = n257 & signy_d3;
  /* fppowtf32.vhdl:6069:7  */
  assign n259 = n256 | n258;
  /* fppowtf32.vhdl:6070:19  */
  assign n260 = infx_d3 & normaly_d3;
  /* fppowtf32.vhdl:6070:40  */
  assign n261 = ~signy_d3;
  /* fppowtf32.vhdl:6070:36  */
  assign n262 = n260 & n261;
  /* fppowtf32.vhdl:6070:7  */
  assign n263 = n259 | n262;
  /* fppowtf32.vhdl:6072:37  */
  assign n264 = oddinty_d1 | eveninty_d1;
  /* fppowtf32.vhdl:6072:20  */
  assign n265 = zerox_d3 & n264;
  /* fppowtf32.vhdl:6072:58  */
  assign n266 = ~signy_d3;
  /* fppowtf32.vhdl:6072:54  */
  assign n267 = n265 & n266;
  /* fppowtf32.vhdl:6073:20  */
  assign n268 = zerox_d3 & infy_d3;
  /* fppowtf32.vhdl:6073:38  */
  assign n269 = ~signy_d3;
  /* fppowtf32.vhdl:6073:34  */
  assign n270 = n268 & n269;
  /* fppowtf32.vhdl:6073:7  */
  assign n271 = n267 | n270;
  /* fppowtf32.vhdl:6074:35  */
  assign n272 = absxltoneandnormal_d3 & infy_d3;
  /* fppowtf32.vhdl:6074:53  */
  assign n273 = ~signy_d3;
  /* fppowtf32.vhdl:6074:49  */
  assign n274 = n272 & n273;
  /* fppowtf32.vhdl:6074:7  */
  assign n275 = n271 | n274;
  /* fppowtf32.vhdl:6075:35  */
  assign n276 = absxgtoneandnormal_d3 & infy_d3;
  /* fppowtf32.vhdl:6075:49  */
  assign n277 = n276 & signy_d3;
  /* fppowtf32.vhdl:6075:7  */
  assign n278 = n275 | n277;
  /* fppowtf32.vhdl:6076:19  */
  assign n279 = infx_d3 & normaly_d3;
  /* fppowtf32.vhdl:6076:36  */
  assign n280 = n279 & signy_d3;
  /* fppowtf32.vhdl:6076:7  */
  assign n281 = n278 | n280;
  /* fppowtf32.vhdl:6079:27  */
  assign n282 = xisoneandnormal & signx;
  /* fppowtf32.vhdl:6079:37  */
  assign n283 = n282 & infy;
  /* fppowtf32.vhdl:6079:7  */
  assign n284 = zeroy | n283;
  /* fppowtf32.vhdl:6080:32  */
  assign n285 = ~signx;
  /* fppowtf32.vhdl:6080:28  */
  assign n286 = xisoneandnormal & n285;
  /* fppowtf32.vhdl:6080:7  */
  assign n287 = n284 | n286;
  /* fppowtf32.vhdl:6081:31  */
  assign n288 = ~zeroy_d2;
  /* fppowtf32.vhdl:6081:27  */
  assign n289 = s_nan_in_d2 & n288;
  /* fppowtf32.vhdl:6081:60  */
  assign n290 = normalx_d2 & signx_d2;
  /* fppowtf32.vhdl:6081:73  */
  assign n291 = n290 & notintnormaly;
  /* fppowtf32.vhdl:6081:45  */
  assign n292 = n289 | n291;
  /* fppowtf32.vhdl:6082:22  */
  assign n293 = signx_d2 & oddinty;
  /* fppowtf32.vhdl:6083:20  */
  assign n295 = {flagsx, 1'b0};
  /* fppowtf32.vhdl:6083:26  */
  assign n296 = {n295, expfieldx};
  /* fppowtf32.vhdl:6083:38  */
  assign n297 = {n296, fracx};
  /* fppowtf32.vhdl:6083:46  */
  assign n299 = {n297, 10'b0000000000};
  /* fppowtf32.vhdl:6084:4  */
  fplogiterative_8_20_0_500_freq500_uid9 fppow_8_10_freq500_uid2log (
    .clk(clk),
    .x(login),
    .r(fppow_8_10_freq500_uid2log_n300));
  /* fppowtf32.vhdl:6088:4  */
  fpmult_8_20_uid62_freq500_uid63 fppow_8_10_freq500_uid2mult (
    .clk(clk),
    .x(lnx),
    .y(Y),
    .r(fppow_8_10_freq500_uid2mult_n303));
  /* fppowtf32.vhdl:6093:4  */
  fpexp_8_10_freq500_uid71 fppow_8_10_freq500_uid2exp (
    .clk(clk),
    .x(p),
    .r(fppow_8_10_freq500_uid2exp_n306));
  /* fppowtf32.vhdl:6097:15  */
  assign n309 = e[20:19]; // extract
  /* fppowtf32.vhdl:6098:40  */
  assign n312 = flagse_d1 == 2'b00;
  /* fppowtf32.vhdl:6098:26  */
  assign n313 = n312 ? 1'b1 : 1'b0;
  /* fppowtf32.vhdl:6099:38  */
  assign n315 = riszerospecialcase_d18 | riszerofromexp;
  /* fppowtf32.vhdl:6100:40  */
  assign n318 = flagse_d1 == 2'b10;
  /* fppowtf32.vhdl:6100:26  */
  assign n319 = n318 ? 1'b1 : 1'b0;
  /* fppowtf32.vhdl:6101:37  */
  assign n321 = risinfspecialcase_d18 | risinffromexp;
  /* fppowtf32.vhdl:6103:17  */
  assign n323 = risnan_d19 ? 2'b11 : n325;
  /* fppowtf32.vhdl:6104:7  */
  assign n325 = riszero ? 2'b00 : n327;
  /* fppowtf32.vhdl:6105:7  */
  assign n327 = risinf ? 2'b10 : 2'b01;
  /* fppowtf32.vhdl:6107:78  */
  assign n330 = risone_d21 ? 18'b011111110000000000 : n331;
  /* fppowtf32.vhdl:6108:17  */
  assign n331 = e_d1[17:0]; // extract
  /* fppowtf32.vhdl:6109:15  */
  assign n332 = {flagr, signr_d19};
  /* fppowtf32.vhdl:6109:27  */
  assign n333 = {n332, r_expfrac};
  /* fppowtf32.vhdl:5885:10  */
  always @(posedge clk)
    n334 <= signx;
  /* fppowtf32.vhdl:5885:10  */
  always @(posedge clk)
    n335 <= signx_d1;
  /* fppowtf32.vhdl:5885:10  */
  always @(posedge clk)
    n336 <= signy;
  /* fppowtf32.vhdl:5885:10  */
  always @(posedge clk)
    n337 <= signy_d1;
  /* fppowtf32.vhdl:5885:10  */
  always @(posedge clk)
    n338 <= signy_d2;
  /* fppowtf32.vhdl:5885:10  */
  always @(posedge clk)
    n339 <= zerox;
  /* fppowtf32.vhdl:5885:10  */
  always @(posedge clk)
    n340 <= zerox_d1;
  /* fppowtf32.vhdl:5885:10  */
  always @(posedge clk)
    n341 <= zerox_d2;
  /* fppowtf32.vhdl:5885:10  */
  always @(posedge clk)
    n342 <= zeroy;
  /* fppowtf32.vhdl:5885:10  */
  always @(posedge clk)
    n343 <= zeroy_d1;
  /* fppowtf32.vhdl:5885:10  */
  always @(posedge clk)
    n344 <= normalx;
  /* fppowtf32.vhdl:5885:10  */
  always @(posedge clk)
    n345 <= normalx_d1;
  /* fppowtf32.vhdl:5885:10  */
  always @(posedge clk)
    n346 <= normaly;
  /* fppowtf32.vhdl:5885:10  */
  always @(posedge clk)
    n347 <= normaly_d1;
  /* fppowtf32.vhdl:5885:10  */
  always @(posedge clk)
    n348 <= normaly_d2;
  /* fppowtf32.vhdl:5885:10  */
  always @(posedge clk)
    n349 <= infx;
  /* fppowtf32.vhdl:5885:10  */
  always @(posedge clk)
    n350 <= infx_d1;
  /* fppowtf32.vhdl:5885:10  */
  always @(posedge clk)
    n351 <= infx_d2;
  /* fppowtf32.vhdl:5885:10  */
  always @(posedge clk)
    n352 <= infy;
  /* fppowtf32.vhdl:5885:10  */
  always @(posedge clk)
    n353 <= infy_d1;
  /* fppowtf32.vhdl:5885:10  */
  always @(posedge clk)
    n354 <= infy_d2;
  /* fppowtf32.vhdl:5885:10  */
  always @(posedge clk)
    n355 <= s_nan_in;
  /* fppowtf32.vhdl:5885:10  */
  always @(posedge clk)
    n356 <= s_nan_in_d1;
  /* fppowtf32.vhdl:5885:10  */
  always @(posedge clk)
    n357 <= absxgtoneandnormal;
  /* fppowtf32.vhdl:5885:10  */
  always @(posedge clk)
    n358 <= absxgtoneandnormal_d1;
  /* fppowtf32.vhdl:5885:10  */
  always @(posedge clk)
    n359 <= absxgtoneandnormal_d2;
  /* fppowtf32.vhdl:5885:10  */
  always @(posedge clk)
    n360 <= absxltoneandnormal;
  /* fppowtf32.vhdl:5885:10  */
  always @(posedge clk)
    n361 <= absxltoneandnormal_d1;
  /* fppowtf32.vhdl:5885:10  */
  always @(posedge clk)
    n362 <= absxltoneandnormal_d2;
  /* fppowtf32.vhdl:5885:10  */
  always @(posedge clk)
    n363 <= z_righty;
  /* fppowtf32.vhdl:5885:10  */
  always @(posedge clk)
    n364 <= weightlsbypre;
  /* fppowtf32.vhdl:5885:10  */
  always @(posedge clk)
    n365 <= weightlsbypre_d1;
  /* fppowtf32.vhdl:5885:10  */
  always @(posedge clk)
    n366 <= oddinty;
  /* fppowtf32.vhdl:5885:10  */
  always @(posedge clk)
    n367 <= eveninty;
  /* fppowtf32.vhdl:5885:10  */
  always @(posedge clk)
    n368 <= risinfspecialcase;
  /* fppowtf32.vhdl:5885:10  */
  always @(posedge clk)
    n369 <= risinfspecialcase_d1;
  /* fppowtf32.vhdl:5885:10  */
  always @(posedge clk)
    n370 <= risinfspecialcase_d2;
  /* fppowtf32.vhdl:5885:10  */
  always @(posedge clk)
    n371 <= risinfspecialcase_d3;
  /* fppowtf32.vhdl:5885:10  */
  always @(posedge clk)
    n372 <= risinfspecialcase_d4;
  /* fppowtf32.vhdl:5885:10  */
  always @(posedge clk)
    n373 <= risinfspecialcase_d5;
  /* fppowtf32.vhdl:5885:10  */
  always @(posedge clk)
    n374 <= risinfspecialcase_d6;
  /* fppowtf32.vhdl:5885:10  */
  always @(posedge clk)
    n375 <= risinfspecialcase_d7;
  /* fppowtf32.vhdl:5885:10  */
  always @(posedge clk)
    n376 <= risinfspecialcase_d8;
  /* fppowtf32.vhdl:5885:10  */
  always @(posedge clk)
    n377 <= risinfspecialcase_d9;
  /* fppowtf32.vhdl:5885:10  */
  always @(posedge clk)
    n378 <= risinfspecialcase_d10;
  /* fppowtf32.vhdl:5885:10  */
  always @(posedge clk)
    n379 <= risinfspecialcase_d11;
  /* fppowtf32.vhdl:5885:10  */
  always @(posedge clk)
    n380 <= risinfspecialcase_d12;
  /* fppowtf32.vhdl:5885:10  */
  always @(posedge clk)
    n381 <= risinfspecialcase_d13;
  /* fppowtf32.vhdl:5885:10  */
  always @(posedge clk)
    n382 <= risinfspecialcase_d14;
  /* fppowtf32.vhdl:5885:10  */
  always @(posedge clk)
    n383 <= risinfspecialcase_d15;
  /* fppowtf32.vhdl:5885:10  */
  always @(posedge clk)
    n384 <= risinfspecialcase_d16;
  /* fppowtf32.vhdl:5885:10  */
  always @(posedge clk)
    n385 <= risinfspecialcase_d17;
  /* fppowtf32.vhdl:5885:10  */
  always @(posedge clk)
    n386 <= riszerospecialcase;
  /* fppowtf32.vhdl:5885:10  */
  always @(posedge clk)
    n387 <= riszerospecialcase_d1;
  /* fppowtf32.vhdl:5885:10  */
  always @(posedge clk)
    n388 <= riszerospecialcase_d2;
  /* fppowtf32.vhdl:5885:10  */
  always @(posedge clk)
    n389 <= riszerospecialcase_d3;
  /* fppowtf32.vhdl:5885:10  */
  always @(posedge clk)
    n390 <= riszerospecialcase_d4;
  /* fppowtf32.vhdl:5885:10  */
  always @(posedge clk)
    n391 <= riszerospecialcase_d5;
  /* fppowtf32.vhdl:5885:10  */
  always @(posedge clk)
    n392 <= riszerospecialcase_d6;
  /* fppowtf32.vhdl:5885:10  */
  always @(posedge clk)
    n393 <= riszerospecialcase_d7;
  /* fppowtf32.vhdl:5885:10  */
  always @(posedge clk)
    n394 <= riszerospecialcase_d8;
  /* fppowtf32.vhdl:5885:10  */
  always @(posedge clk)
    n395 <= riszerospecialcase_d9;
  /* fppowtf32.vhdl:5885:10  */
  always @(posedge clk)
    n396 <= riszerospecialcase_d10;
  /* fppowtf32.vhdl:5885:10  */
  always @(posedge clk)
    n397 <= riszerospecialcase_d11;
  /* fppowtf32.vhdl:5885:10  */
  always @(posedge clk)
    n398 <= riszerospecialcase_d12;
  /* fppowtf32.vhdl:5885:10  */
  always @(posedge clk)
    n399 <= riszerospecialcase_d13;
  /* fppowtf32.vhdl:5885:10  */
  always @(posedge clk)
    n400 <= riszerospecialcase_d14;
  /* fppowtf32.vhdl:5885:10  */
  always @(posedge clk)
    n401 <= riszerospecialcase_d15;
  /* fppowtf32.vhdl:5885:10  */
  always @(posedge clk)
    n402 <= riszerospecialcase_d16;
  /* fppowtf32.vhdl:5885:10  */
  always @(posedge clk)
    n403 <= riszerospecialcase_d17;
  /* fppowtf32.vhdl:5885:10  */
  always @(posedge clk)
    n404 <= risone;
  /* fppowtf32.vhdl:5885:10  */
  always @(posedge clk)
    n405 <= risone_d1;
  /* fppowtf32.vhdl:5885:10  */
  always @(posedge clk)
    n406 <= risone_d2;
  /* fppowtf32.vhdl:5885:10  */
  always @(posedge clk)
    n407 <= risone_d3;
  /* fppowtf32.vhdl:5885:10  */
  always @(posedge clk)
    n408 <= risone_d4;
  /* fppowtf32.vhdl:5885:10  */
  always @(posedge clk)
    n409 <= risone_d5;
  /* fppowtf32.vhdl:5885:10  */
  always @(posedge clk)
    n410 <= risone_d6;
  /* fppowtf32.vhdl:5885:10  */
  always @(posedge clk)
    n411 <= risone_d7;
  /* fppowtf32.vhdl:5885:10  */
  always @(posedge clk)
    n412 <= risone_d8;
  /* fppowtf32.vhdl:5885:10  */
  always @(posedge clk)
    n413 <= risone_d9;
  /* fppowtf32.vhdl:5885:10  */
  always @(posedge clk)
    n414 <= risone_d10;
  /* fppowtf32.vhdl:5885:10  */
  always @(posedge clk)
    n415 <= risone_d11;
  /* fppowtf32.vhdl:5885:10  */
  always @(posedge clk)
    n416 <= risone_d12;
  /* fppowtf32.vhdl:5885:10  */
  always @(posedge clk)
    n417 <= risone_d13;
  /* fppowtf32.vhdl:5885:10  */
  always @(posedge clk)
    n418 <= risone_d14;
  /* fppowtf32.vhdl:5885:10  */
  always @(posedge clk)
    n419 <= risone_d15;
  /* fppowtf32.vhdl:5885:10  */
  always @(posedge clk)
    n420 <= risone_d16;
  /* fppowtf32.vhdl:5885:10  */
  always @(posedge clk)
    n421 <= risone_d17;
  /* fppowtf32.vhdl:5885:10  */
  always @(posedge clk)
    n422 <= risone_d18;
  /* fppowtf32.vhdl:5885:10  */
  always @(posedge clk)
    n423 <= risone_d19;
  /* fppowtf32.vhdl:5885:10  */
  always @(posedge clk)
    n424 <= risone_d20;
  /* fppowtf32.vhdl:5885:10  */
  always @(posedge clk)
    n425 <= risnan;
  /* fppowtf32.vhdl:5885:10  */
  always @(posedge clk)
    n426 <= risnan_d1;
  /* fppowtf32.vhdl:5885:10  */
  always @(posedge clk)
    n427 <= risnan_d2;
  /* fppowtf32.vhdl:5885:10  */
  always @(posedge clk)
    n428 <= risnan_d3;
  /* fppowtf32.vhdl:5885:10  */
  always @(posedge clk)
    n429 <= risnan_d4;
  /* fppowtf32.vhdl:5885:10  */
  always @(posedge clk)
    n430 <= risnan_d5;
  /* fppowtf32.vhdl:5885:10  */
  always @(posedge clk)
    n431 <= risnan_d6;
  /* fppowtf32.vhdl:5885:10  */
  always @(posedge clk)
    n432 <= risnan_d7;
  /* fppowtf32.vhdl:5885:10  */
  always @(posedge clk)
    n433 <= risnan_d8;
  /* fppowtf32.vhdl:5885:10  */
  always @(posedge clk)
    n434 <= risnan_d9;
  /* fppowtf32.vhdl:5885:10  */
  always @(posedge clk)
    n435 <= risnan_d10;
  /* fppowtf32.vhdl:5885:10  */
  always @(posedge clk)
    n436 <= risnan_d11;
  /* fppowtf32.vhdl:5885:10  */
  always @(posedge clk)
    n437 <= risnan_d12;
  /* fppowtf32.vhdl:5885:10  */
  always @(posedge clk)
    n438 <= risnan_d13;
  /* fppowtf32.vhdl:5885:10  */
  always @(posedge clk)
    n439 <= risnan_d14;
  /* fppowtf32.vhdl:5885:10  */
  always @(posedge clk)
    n440 <= risnan_d15;
  /* fppowtf32.vhdl:5885:10  */
  always @(posedge clk)
    n441 <= risnan_d16;
  /* fppowtf32.vhdl:5885:10  */
  always @(posedge clk)
    n442 <= risnan_d17;
  /* fppowtf32.vhdl:5885:10  */
  always @(posedge clk)
    n443 <= risnan_d18;
  /* fppowtf32.vhdl:5885:10  */
  always @(posedge clk)
    n444 <= signr;
  /* fppowtf32.vhdl:5885:10  */
  always @(posedge clk)
    n445 <= signr_d1;
  /* fppowtf32.vhdl:5885:10  */
  always @(posedge clk)
    n446 <= signr_d2;
  /* fppowtf32.vhdl:5885:10  */
  always @(posedge clk)
    n447 <= signr_d3;
  /* fppowtf32.vhdl:5885:10  */
  always @(posedge clk)
    n448 <= signr_d4;
  /* fppowtf32.vhdl:5885:10  */
  always @(posedge clk)
    n449 <= signr_d5;
  /* fppowtf32.vhdl:5885:10  */
  always @(posedge clk)
    n450 <= signr_d6;
  /* fppowtf32.vhdl:5885:10  */
  always @(posedge clk)
    n451 <= signr_d7;
  /* fppowtf32.vhdl:5885:10  */
  always @(posedge clk)
    n452 <= signr_d8;
  /* fppowtf32.vhdl:5885:10  */
  always @(posedge clk)
    n453 <= signr_d9;
  /* fppowtf32.vhdl:5885:10  */
  always @(posedge clk)
    n454 <= signr_d10;
  /* fppowtf32.vhdl:5885:10  */
  always @(posedge clk)
    n455 <= signr_d11;
  /* fppowtf32.vhdl:5885:10  */
  always @(posedge clk)
    n456 <= signr_d12;
  /* fppowtf32.vhdl:5885:10  */
  always @(posedge clk)
    n457 <= signr_d13;
  /* fppowtf32.vhdl:5885:10  */
  always @(posedge clk)
    n458 <= signr_d14;
  /* fppowtf32.vhdl:5885:10  */
  always @(posedge clk)
    n459 <= signr_d15;
  /* fppowtf32.vhdl:5885:10  */
  always @(posedge clk)
    n460 <= signr_d16;
  /* fppowtf32.vhdl:5885:10  */
  always @(posedge clk)
    n461 <= signr_d17;
  /* fppowtf32.vhdl:5885:10  */
  always @(posedge clk)
    n462 <= signr_d18;
  /* fppowtf32.vhdl:5885:10  */
  always @(posedge clk)
    n463 <= e;
  /* fppowtf32.vhdl:5885:10  */
  always @(posedge clk)
    n464 <= flagse;
endmodule

